VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Onchip_RCO
  CLASS BLOCK ;
  FOREIGN tt_um_Onchip_RCO ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[2]
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 2.100000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNAGATEAREA 15.400000 ;
    ANTENNADIFFAREA 24.855999 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  PIN ua[1]
    ANTENNADIFFAREA 1.800000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN vss
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT 120.605 31.920 120.615 31.930 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.440 31.890 136.450 31.900 ;
    END
    PORT
      LAYER met1 ;
        RECT 123.030 20.205 123.040 20.215 ;
    END
    PORT
      LAYER met1 ;
        RECT 125.625 20.205 125.635 20.215 ;
    END
    PORT
      LAYER met1 ;
        RECT 127.575 20.205 127.585 20.215 ;
    END
    PORT
      LAYER met1 ;
        RECT 129.525 20.205 129.535 20.215 ;
    END
    PORT
      LAYER met1 ;
        RECT 131.475 20.205 131.485 20.215 ;
    END
    PORT
      LAYER met1 ;
        RECT 123.855 20.205 123.865 20.215 ;
    END
    PORT
      LAYER met1 ;
        RECT 125.805 20.205 125.815 20.215 ;
    END
    PORT
      LAYER met1 ;
        RECT 127.755 20.205 127.765 20.215 ;
    END
    PORT
      LAYER met1 ;
        RECT 129.705 20.205 129.715 20.215 ;
    END
    PORT
      LAYER met1 ;
        RECT 131.655 20.205 131.665 20.215 ;
    END
    PORT
      LAYER met1 ;
        RECT 133.605 20.205 133.615 20.215 ;
    END
    PORT
      LAYER met1 ;
        RECT 133.425 20.205 133.435 20.215 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.355 21.735 123.365 21.745 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.595 21.735 125.605 21.745 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.545 21.735 127.555 21.745 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.495 21.735 129.505 21.745 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.445 21.735 131.455 21.745 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.885 18.675 123.895 18.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.835 18.675 125.845 18.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.785 18.675 127.795 18.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.735 18.675 129.745 18.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.685 18.675 131.695 18.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.635 18.675 133.645 18.685 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.395 21.735 133.405 21.745 ;
    END
  END vss
  PIN out
    ANTENNADIFFAREA 1.800000 ;
    PORT
      LAYER met1 ;
        RECT 136.635 25.930 136.645 25.940 ;
    END
    PORT
      LAYER met1 ;
        RECT 127.510 25.110 127.520 25.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 129.460 25.110 129.470 25.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 131.410 25.110 131.420 25.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 123.920 15.300 123.930 15.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 125.870 15.300 125.880 15.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 127.820 15.300 127.830 15.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 129.770 15.300 129.780 15.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 131.720 15.300 131.730 15.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 133.670 15.300 133.680 15.310 ;
    END
    PORT
      LAYER met1 ;
        RECT 133.360 25.110 133.370 25.120 ;
    END
    PORT
      LAYER met1 ;
        RECT 125.560 25.110 125.570 25.120 ;
    END
  END out
  PIN vrst
    ANTENNAGATEAREA 2.100000 ;
    PORT
      LAYER met1 ;
        RECT 122.440 24.310 122.450 24.320 ;
    END
  END vrst
  PIN vdd
    ANTENNAGATEAREA 15.400000 ;
    ANTENNADIFFAREA 24.855999 ;
    PORT
      LAYER met1 ;
        RECT 123.035 31.985 123.045 31.995 ;
    END
    PORT
      LAYER met1 ;
        RECT 125.665 31.985 125.675 31.995 ;
    END
    PORT
      LAYER met1 ;
        RECT 127.615 31.985 127.625 31.995 ;
    END
    PORT
      LAYER met1 ;
        RECT 129.565 31.985 129.575 31.995 ;
    END
    PORT
      LAYER met1 ;
        RECT 131.515 31.985 131.525 31.995 ;
    END
    PORT
      LAYER met1 ;
        RECT 123.815 8.425 123.825 8.435 ;
    END
    PORT
      LAYER met1 ;
        RECT 125.765 8.425 125.775 8.435 ;
    END
    PORT
      LAYER met1 ;
        RECT 127.715 8.425 127.725 8.435 ;
    END
    PORT
      LAYER met1 ;
        RECT 129.665 8.425 129.675 8.435 ;
    END
    PORT
      LAYER met1 ;
        RECT 131.615 8.425 131.625 8.435 ;
    END
    PORT
      LAYER met1 ;
        RECT 133.565 8.425 133.575 8.435 ;
    END
    PORT
      LAYER met1 ;
        RECT 133.465 31.985 133.475 31.995 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.390 29.955 123.400 29.965 ;
    END
  END vdd
  PIN in
    ANTENNAGATEAREA 1.050000 ;
    ANTENNADIFFAREA 0.900000 ;
    PORT
      LAYER met1 ;
        RECT 125.765 25.095 125.775 25.105 ;
    END
    PORT
      LAYER met1 ;
        RECT 127.715 25.095 127.725 25.105 ;
    END
    PORT
      LAYER met1 ;
        RECT 129.665 25.095 129.675 25.105 ;
    END
    PORT
      LAYER met1 ;
        RECT 125.665 15.315 125.675 15.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 127.615 15.315 127.625 15.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 129.565 15.315 129.575 15.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 131.515 15.315 131.525 15.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 133.465 15.315 133.475 15.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 135.415 15.315 135.425 15.325 ;
    END
    PORT
      LAYER met1 ;
        RECT 131.615 25.095 131.625 25.105 ;
    END
    PORT
      LAYER met1 ;
        RECT 123.815 25.095 123.825 25.105 ;
    END
  END in
  PIN vctrn
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER met3 ;
        RECT 122.425 19.540 122.435 19.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 122.425 20.870 122.435 20.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.640 20.870 125.650 20.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.590 20.870 127.600 20.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.540 20.870 129.550 20.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.490 20.870 131.500 20.880 ;
    END
    PORT
      LAYER met3 ;
        RECT 123.840 19.540 123.850 19.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.790 19.540 125.800 19.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.740 19.540 127.750 19.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.690 19.540 129.700 19.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.640 19.540 131.650 19.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.590 19.540 133.600 19.550 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.440 20.870 133.450 20.880 ;
    END
  END vctrn
  PIN vctrp
    ANTENNAGATEAREA 8.400000 ;
    ANTENNADIFFAREA 0.900000 ;
    PORT
      LAYER met3 ;
        RECT 123.845 9.045 123.855 9.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 125.795 9.045 125.805 9.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 127.745 9.045 127.755 9.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 129.695 9.045 129.705 9.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 131.645 9.045 131.655 9.055 ;
    END
    PORT
      LAYER met3 ;
        RECT 133.595 9.045 133.605 9.055 ;
    END
  END vctrp
  OBS
      LAYER nwell ;
        RECT 122.665 8.050 136.345 32.370 ;
      LAYER li1 ;
        RECT 122.940 8.230 135.975 32.190 ;
      LAYER met1 ;
        RECT 120.425 31.705 122.755 32.190 ;
        RECT 123.325 31.705 125.385 32.190 ;
        RECT 125.955 31.705 127.335 32.190 ;
        RECT 127.905 31.705 129.285 32.190 ;
        RECT 129.855 31.705 131.235 32.190 ;
        RECT 131.805 31.705 133.185 32.190 ;
        RECT 133.755 31.705 138.760 32.190 ;
        RECT 120.425 26.220 138.760 31.705 ;
        RECT 120.425 25.650 136.355 26.220 ;
        RECT 136.925 25.650 138.760 26.220 ;
        RECT 120.425 25.400 138.760 25.650 ;
        RECT 120.425 25.385 125.280 25.400 ;
        RECT 125.850 25.385 127.230 25.400 ;
        RECT 127.800 25.385 129.180 25.400 ;
        RECT 129.750 25.385 131.130 25.400 ;
        RECT 131.700 25.385 133.080 25.400 ;
        RECT 120.425 24.815 123.535 25.385 ;
        RECT 124.105 24.830 125.280 25.385 ;
        RECT 126.055 24.830 127.230 25.385 ;
        RECT 128.005 24.830 129.180 25.385 ;
        RECT 129.955 24.830 131.130 25.385 ;
        RECT 131.905 24.830 133.080 25.385 ;
        RECT 133.650 24.830 138.760 25.400 ;
        RECT 124.105 24.815 125.485 24.830 ;
        RECT 126.055 24.815 127.435 24.830 ;
        RECT 128.005 24.815 129.385 24.830 ;
        RECT 129.955 24.815 131.335 24.830 ;
        RECT 131.905 24.815 138.760 24.830 ;
        RECT 120.425 24.600 138.760 24.815 ;
        RECT 120.425 24.030 122.160 24.600 ;
        RECT 122.730 24.030 138.760 24.600 ;
        RECT 120.425 20.495 138.760 24.030 ;
        RECT 120.425 19.925 122.750 20.495 ;
        RECT 123.320 19.925 123.575 20.495 ;
        RECT 124.145 19.925 125.345 20.495 ;
        RECT 126.095 19.925 127.295 20.495 ;
        RECT 128.045 19.925 129.245 20.495 ;
        RECT 129.995 19.925 131.195 20.495 ;
        RECT 131.945 19.925 133.145 20.495 ;
        RECT 133.895 19.925 138.760 20.495 ;
        RECT 120.425 15.605 138.760 19.925 ;
        RECT 120.425 15.590 125.385 15.605 ;
        RECT 125.955 15.590 127.335 15.605 ;
        RECT 127.905 15.590 129.285 15.605 ;
        RECT 129.855 15.590 131.235 15.605 ;
        RECT 131.805 15.590 133.185 15.605 ;
        RECT 133.755 15.590 135.135 15.605 ;
        RECT 120.425 15.020 123.640 15.590 ;
        RECT 124.210 15.035 125.385 15.590 ;
        RECT 126.160 15.035 127.335 15.590 ;
        RECT 128.110 15.035 129.285 15.590 ;
        RECT 130.060 15.035 131.235 15.590 ;
        RECT 132.010 15.035 133.185 15.590 ;
        RECT 133.960 15.035 135.135 15.590 ;
        RECT 135.705 15.035 138.760 15.605 ;
        RECT 124.210 15.020 125.590 15.035 ;
        RECT 126.160 15.020 127.540 15.035 ;
        RECT 128.110 15.020 129.490 15.035 ;
        RECT 130.060 15.020 131.440 15.035 ;
        RECT 132.010 15.020 133.390 15.035 ;
        RECT 133.960 15.020 138.760 15.035 ;
        RECT 120.425 8.715 138.760 15.020 ;
        RECT 120.425 8.230 123.535 8.715 ;
        RECT 124.105 8.230 125.485 8.715 ;
        RECT 126.055 8.230 127.435 8.715 ;
        RECT 128.005 8.230 129.385 8.715 ;
        RECT 129.955 8.230 131.335 8.715 ;
        RECT 131.905 8.230 133.285 8.715 ;
        RECT 133.855 8.230 138.760 8.715 ;
      LAYER met2 ;
        RECT 120.425 8.230 138.760 32.190 ;
      LAYER met3 ;
        RECT 1.000 30.365 141.145 41.895 ;
        RECT 1.000 29.555 122.990 30.365 ;
        RECT 123.800 29.555 141.145 30.365 ;
        RECT 1.000 22.145 141.145 29.555 ;
        RECT 1.000 21.335 122.955 22.145 ;
        RECT 123.765 21.335 125.195 22.145 ;
        RECT 126.005 21.335 127.145 22.145 ;
        RECT 127.955 21.335 129.095 22.145 ;
        RECT 129.905 21.335 131.045 22.145 ;
        RECT 131.855 21.335 132.995 22.145 ;
        RECT 133.805 21.335 141.145 22.145 ;
        RECT 1.000 21.280 141.145 21.335 ;
        RECT 1.000 20.470 122.025 21.280 ;
        RECT 122.835 20.470 125.240 21.280 ;
        RECT 126.050 20.470 127.190 21.280 ;
        RECT 128.000 20.470 129.140 21.280 ;
        RECT 129.950 20.470 131.090 21.280 ;
        RECT 131.900 20.470 133.040 21.280 ;
        RECT 133.850 20.470 141.145 21.280 ;
        RECT 1.000 19.950 141.145 20.470 ;
        RECT 1.000 19.140 122.025 19.950 ;
        RECT 122.835 19.140 123.440 19.950 ;
        RECT 124.250 19.140 125.390 19.950 ;
        RECT 126.200 19.140 127.340 19.950 ;
        RECT 128.150 19.140 129.290 19.950 ;
        RECT 130.100 19.140 131.240 19.950 ;
        RECT 132.050 19.140 133.190 19.950 ;
        RECT 134.000 19.140 141.145 19.950 ;
        RECT 1.000 19.085 141.145 19.140 ;
        RECT 1.000 18.275 123.485 19.085 ;
        RECT 124.295 18.275 125.435 19.085 ;
        RECT 126.245 18.275 127.385 19.085 ;
        RECT 128.195 18.275 129.335 19.085 ;
        RECT 130.145 18.275 131.285 19.085 ;
        RECT 132.095 18.275 133.235 19.085 ;
        RECT 134.045 18.275 141.145 19.085 ;
        RECT 1.000 9.455 141.145 18.275 ;
        RECT 1.000 8.645 123.445 9.455 ;
        RECT 124.255 8.645 125.395 9.455 ;
        RECT 126.205 8.645 127.345 9.455 ;
        RECT 128.155 8.645 129.295 9.455 ;
        RECT 130.105 8.645 131.245 9.455 ;
        RECT 132.055 8.645 133.195 9.455 ;
        RECT 134.005 8.645 141.145 9.455 ;
        RECT 1.000 8.230 141.145 8.645 ;
      LAYER met4 ;
        RECT 6.000 224.360 30.270 224.760 ;
        RECT 31.370 224.360 33.030 224.760 ;
        RECT 34.130 224.360 35.790 224.760 ;
        RECT 36.890 224.360 38.550 224.760 ;
        RECT 39.650 224.360 41.310 224.760 ;
        RECT 42.410 224.360 44.070 224.760 ;
        RECT 45.170 224.360 46.830 224.760 ;
        RECT 47.930 224.360 49.590 224.760 ;
        RECT 50.690 224.360 52.350 224.760 ;
        RECT 53.450 224.360 55.110 224.760 ;
        RECT 56.210 224.360 57.870 224.760 ;
        RECT 58.970 224.360 60.630 224.760 ;
        RECT 61.730 224.360 63.390 224.760 ;
        RECT 64.490 224.360 66.150 224.760 ;
        RECT 67.250 224.360 68.910 224.760 ;
        RECT 70.010 224.360 71.670 224.760 ;
        RECT 72.770 224.360 74.430 224.760 ;
        RECT 75.530 224.360 77.190 224.760 ;
        RECT 78.290 224.360 79.950 224.760 ;
        RECT 81.050 224.360 82.710 224.760 ;
        RECT 83.810 224.360 85.470 224.760 ;
        RECT 86.570 224.360 88.230 224.760 ;
        RECT 89.330 224.360 90.990 224.760 ;
        RECT 92.090 224.360 93.750 224.760 ;
        RECT 94.850 224.360 96.510 224.760 ;
        RECT 97.610 224.360 99.270 224.760 ;
        RECT 100.370 224.360 102.030 224.760 ;
        RECT 103.130 224.360 104.790 224.760 ;
        RECT 105.890 224.360 107.550 224.760 ;
        RECT 108.650 224.360 110.310 224.760 ;
        RECT 111.410 224.360 113.070 224.760 ;
        RECT 114.170 224.360 115.830 224.760 ;
        RECT 116.930 224.360 118.590 224.760 ;
        RECT 119.690 224.360 121.350 224.760 ;
        RECT 122.450 224.360 124.110 224.760 ;
        RECT 125.210 224.360 126.870 224.760 ;
        RECT 127.970 224.360 129.630 224.760 ;
        RECT 130.730 224.360 132.390 224.760 ;
        RECT 133.490 224.360 135.150 224.760 ;
        RECT 136.250 224.360 137.910 224.760 ;
        RECT 139.010 224.360 140.670 224.760 ;
        RECT 141.770 224.360 143.430 224.760 ;
        RECT 144.530 224.360 146.190 224.760 ;
        RECT 147.290 224.360 152.715 224.760 ;
        RECT 6.000 221.160 152.715 224.360 ;
        RECT 6.400 32.330 152.715 221.160 ;
        RECT 6.400 31.520 120.205 32.330 ;
        RECT 121.015 32.300 152.715 32.330 ;
        RECT 121.015 31.520 136.040 32.300 ;
        RECT 6.400 31.490 136.040 31.520 ;
        RECT 136.850 31.490 152.715 32.300 ;
        RECT 6.400 4.600 152.715 31.490 ;
        RECT 6.000 1.400 152.715 4.600 ;
        RECT 6.000 0.000 16.170 1.400 ;
        RECT 17.870 0.000 35.490 1.400 ;
        RECT 37.190 0.000 54.810 1.400 ;
        RECT 56.510 0.000 74.130 1.400 ;
        RECT 75.830 0.000 93.450 1.400 ;
        RECT 95.150 0.000 112.770 1.400 ;
        RECT 114.470 0.000 132.090 1.400 ;
        RECT 133.790 0.000 151.410 1.400 ;
  END
END tt_um_Onchip_RCO
END LIBRARY

