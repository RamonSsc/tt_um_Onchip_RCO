magic
tech sky130a
timestamp 1762644065
<< checkpaint >>
rect 0 0 2 1
<< l70d20 >>
rect 0 0 2 1
<< l71d20 >>
rect 0 0 2 1
<< end >>
