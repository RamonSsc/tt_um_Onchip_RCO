  X �  	    �  	     LIB  >A�7KƧ�9D�/��ZT �  	    �  	     tt_um_Onchip_RCO    F   , �  d� �  f:   f:   d� �  d�      F   , ��  �� ��  �� ��  �� ��  �� ��  ��      F   , �  �� �  �x �  �x �  �� �  ��      F   , 	  �� 	  �x �  �x �  �� 	  ��      F   , �/  �� �/  ��    ��    �� �/  ��      F   , �.  �� �.  �x �  �x �  �� �.  ��      F   , k  �� k  �� S  �� S  �� k  ��      F   , �U  �� �U  �x �=  �x �=  �� �U  ��      F   , ��  �� ��  �x �y  �x �y  �� ��  ��      F   , ��  �� ��  �� ��  �� ��  �� ��  ��      F   ,  �  ��  �  �x  p  �x  p  ��  �  ��      F   ,  �  ��  �  ��  �  ��  �  ��  �  ��      F   , �a  S\ �a  V| �=  V| �=  S\ �a  S\      F   , #�  K� #�  M 'Y  M 'Y  K� #�  K�      F   , #�  P� #�  RD 'Y  RD 'Y  P� #�  P�   	   F   !     �  �o  u �_  u   	   F   !     �  �  u ��  u   	   F   !     �  �  u ��  u   	   F   !     �  ��  (� ��  (�   	   F   !     �  �_  (� �o  (�   	   F   !     �  ��  (� �  (�   	   F   !     �  ��  (� �  (�   	   F   !     �  9  (� 
I  (�   	   F   !     �  �  (� �  (�   	   F   !     �  
I  u 9  u   	   F   !     �  ��  u ��  u   	   F   !     J  �  z] �  z]   	   F   !     J  �  z] �T  z]   	   F   !     J  �T  z] �  z]   	   F   !     J  �  #� �z  #�   	   F   !     J  �  #� �  #�   	   F   !     J  �T  #� �  #�   	   F   !     J  �  #� �T  #�   	   F   !     J  	�  #� �  #�   	   F   !     J  .  #� 	�  #�   	   F   !     J  �  z] 	�  z]   	   F   !     J  �z  z] �  z]   	   F   !     �  �_  T� �o  T�   	   F   !     �  ��  T� �  T�   	   F   !     �  ��  T� �  T�   	   F   !     �  ��  H� ��  H�   	   F   !     �  �o  H� �_  H�   	   F   !     �  �  H� ��  H�   	   F   !     �  �  H� ��  H�   	   F   !     �  
I  H� 9  H�   	   F   !     �  �  H� �  H�   	   F   !     �  9  T� 
I  T�   	   F   !     �  ��  T� ��  T�   	   F   !     J  �  Q� �  Q�   	   F   !     J  �  Q� �T  Q�   	   F   !     J  �T  Q� �  Q�   	   F   !     J  �  LY �z  LY   	   F   !     J  �  LY �  LY   	   F   !     J  �T  LY �  LY   	   F   !     J  �  LY �T  LY   	   F   !     J  	�  LY �  LY   	   F   !     J  .  LY 	�  LY   	   F   !     J  �  Q� 	�  Q�   	   F   !     J  �z  Q� �  Q�   	   F   !     �  �z  T� ��  T�   	   F   !     J  'Y  Q� ��  Q�   	   F   !     �  �  T� �P  T�   	   F   !     �  �  u �P  u   	   F   !     �  �  (� �)  (�   	   F   !     J  �  z] �P  z]   	   F   !     J  �P  z] �i  z]   	   F   !     J  �  #� �i  #�   	   F   !     J  �P  Q� ֛  Q�   	   F   !     J  �z  LY �  LY   	   F   !     J  ٧  T �a  T   	   F   !     J  'Y  LY ��  LY   	   F   !     �   �  �� �  ��   	   F   !     �   �  �� �  ��      F   , ��  S� ��  U� �y  U� �y  S� ��  S�      F   , ��  G� ��  I� �y  I� �y  G� ��  G�      F   , �  N* �  O� �  O� �  N* �  N*      F   , ��  N* ��  O� �y  O� �y  N* ��  N*      F   , �U  N* �U  O� �=  O� �=  N* �U  N*      F   , �  G� �  I� ��  I� ��  G� �  G�      F   , �  '� �  )� ��  )� ��  '� �  '�      F   , k  t k  v S  v S  t k  t      F   , �/  t �/  v    v    t �/  t      F   , k  |. k  }� S  }� S  |. k  |.      F   , k  |. k  }� S  }� S  |. k  |.      F   , �/  |. �/  }�    }�    |. �/  |.      F   , �/  |. �/  }�    }�    |. �/  |.      F   ,   W   X\ �  X\ �  W   W      F   , ��  P� ��  R0 �>  R0 �>  P� ��  P�      F   , �j  P� �j  R0 ��  R0 ��  P� �j  P�      F   ,   P�   R0 z  R0 z  P�   P�      F   , ��  y� ��  { �>  { �>  y� ��  y�      F   , �j  y� �j  { ��  { ��  y� �j  y�      F   ,   y�   { z  { z  y�   y�      F   , ��  S� ��  U� �  U� �  S� ��  S�      F   , 9  S� 9  U� �  U� �  S� 9  S�      F   , �  S� �  U� 
I  U� 
I  S� �  S�      F   , ��  t ��  v �  v �  t ��  t      F   , 9  t 9  v �  v �  t 9  t      F   , �  t �  v 
I  v 
I  t �  t      F   , ��  t ��  v �  v �  t ��  t      F   , 9  t 9  v �  v �  t 9  t      F   , �  S� �  U� ��  U� ��  S� �  S�      F   , ��  S� ��  U�  !  U�  !  S� ��  S�      F   , �  S� �  U� �  U� �  S� �  S�      F   , M  S� M  U� �  U� �  S� M  S�      F   , ��  S� ��  U� �  U� �  S� ��  S�      F   , 9  S� 9  U� �  U� �  S� 9  S�      F   , �  t �  v ��  v ��  t �  t      F   , ��  t ��  v  !  v  !  t ��  t      F   , k  p! k  qk S  qk S  p! k  p!      F   , M  t M  v �  v �  t M  t      F   , �_  S� �_  U� ��  U� ��  S� �_  S�      F   , ��  t ��  v �o  v �o  t ��  t      F   , �5  S\ �5  T� ٧  T� ٧  S\ �5  S\      F   , �.  P� �.  R0 �  R0 �  P� �.  P�      F   , �i  y� �i  { ��  { ��  y� �i  y�      F   , �_  t �_  v ��  v ��  t �_  t      F   , �_  t �_  v ��  v ��  t �_  t      F   , ��  t ��  v �o  v �o  t ��  t      F   , �(  P� �(  R0 �  R0 �  P� �(  P�      F   , ��  t ��  v ��  v ��  t ��  t      F   , ��  t ��  v �3  v �3  t ��  t      F   , �s  S� �s  U� ��  U� ��  S� �s  S�      F   , �  P� �  R0 �  R0 �  P� �  P�      F   , �.  y� �.  { �  { �  y� �.  y�      F   , �U  S� �U  U� �=  U� �=  S� �U  S�      F   , �  P� �  R0 �s  R0 �s  P� �  P�      F   , ��  S� ��  U� �G  U� �G  S� ��  S�      F   , �_  S� �_  U� ��  U� ��  S� �_  S�      F   , ��  S� ��  U� �o  U� �o  S� ��  S�      F   , ��  |. ��  }� ��  }� ��  |. ��  |.      F   , �  y� �  { �  { �  y� �  y�      F   , ��  S� ��  U� �3  U� �3  S� ��  S�      F   , �s  t �s  v ��  v ��  t �s  t      F   , ��  S� ��  U� �o  U� �o  S� ��  S�      F   , ��  |. ��  }� ��  }� ��  |. ��  |.      F   , ��  |. ��  }� ��  }� ��  |. ��  |.      F   , ��  |. ��  }� ��  }� ��  |. ��  |.      F   , ��  t ��  v �G  v �G  t ��  t      F   , �  P� �  R0 �  R0 �  P� �  P�      F   , �.  P� �.  R0 �  R0 �  P� �.  P�      F   , �P  y� �P  { ��  { ��  y� �P  y�      F   , �U  G� �U  I� �=  I� �=  G� �U  G�      F   , �  K� �  L� �  L� �  K� �  K�      F   , ��  G� ��  I� �3  I� �3  G� ��  G�      F   , �_  G� �_  I� ��  I� ��  G� �_  G�      F   , �K  G� �K  I� �  I� �  G� �K  G�      F   , ��  G� ��  I� �[  I� �[  G� ��  G�      F   , ��  G� ��  I� �o  I� �o  G� ��  G�      F   , �.  K� �.  L� �  L� �  K� �.  K�      F   , �i  "� �i  $, ��  $, ��  "� �i  "�      F   , ��   & ��  !� ��  !� ��   & ��   &      F   , ��   & ��  !� ��  !� ��   & ��   &      F   , ��   & ��  !� ��  !� ��   & ��   &      F   , �_  G� �_  I� ��  I� ��  G� �_  G�      F   , ��  G� ��  I� �o  I� �o  G� ��  G�      F   , ��  '� ��  )� �3  )� �3  '� ��  '�      F   , �_  '� �_  )� ��  )� ��  '� �_  '�      F   , ��  '� ��  )� �o  )� �o  '� ��  '�      F   , ��   & ��  !� ��  !� ��   & ��   &      F   , �  "� �  $, �  $, �  "� �  "�      F   , �K  '� �K  )� �  )� �  '� �K  '�      F   , ��  '� ��  )� �[  )� �[  '� ��  '�      F   , �.  "� �.  $, �  $, �  "� �.  "�      F   , �  K� �  L� �s  L� �s  K� �  K�      F   , ��  '� ��  )� ��  )� ��  '� ��  '�      F   , �_  '� �_  )� ��  )� ��  '� �_  '�      F   , ��  '� ��  )� �o  )� �o  '� ��  '�      F   , ��  '� ��  )� ��  )� ��  '� ��  '�      F   , k   & k  !� S  !� S   & k   &      F   , k   & k  !� S  !� S   & k   &      F   , �/   & �/  !�    !�     & �/   &      F   , ��  "� ��  $, �>  $, �>  "� ��  "�      F   , �j  "� �j  $, ��  $, ��  "� �j  "�      F   , �%  G� �%  I� ��  I� ��  G� �%  G�      F   , �  G� �  I� 5  I� 5  G� �  G�      F   , a  G� a  I� �  I� �  G� a  G�      F   ,   "�   $, z  $, z  "�   "�      F   , �  "� �  $,   $,   "� �  "�      F   , ��  K� ��  L� �>  L� �>  K� ��  K�      F   , ��  '� ��  )� �  )� �  '� ��  '�      F   , 9  '� 9  )� �  )� �  '� 9  '�      F   , �  '� �  )� 
I  )� 
I  '� �  '�      F   , �j  K� �j  L� ��  L� ��  K� �j  K�      F   , ��  G� ��  I� �  I� �  G� ��  G�      F   , 9  G� 9  I� �  I� �  G� 9  G�      F   , �  G� �  I� 
I  I� 
I  G� �  G�      F   , u  G� u  I� �  I� �  G� u  G�      F   ,   K�   L� z  L� z  K�   K�      F   , �  K� �  L�   L�   K� �  K�      F   , �/   & �/  !�    !�     & �/   &      F   , k  '� k  )� S  )� S  '� k  '�      F   , �  G� �  I� �  I� �  G� �  G�      F   , �/  '� �/  )�    )�    '� �/  '�      F   , ��  '� ��  )� �  )� �  '� ��  '�      F   , 9  '� 9  )� �  )� �  '� 9  '�      F   , �%  '� �%  )� ��  )� ��  '� �%  '�      F   , �  '� �  )� 5  )� 5  '� �  '�      F   , a  '� a  )� �  )� �  '� a  '�      F   , �  '� �  )� 
I  )� 
I  '� �  '�      F   , u  '� u  )� �  )� �  '� u  '�      F   , ��  G� ��  I� �  I� �  G� ��  G�      F   , 9  G� 9  I� �  I� �  G� 9  G�      F   , �  G� �  I� 
I  I� 
I  G� �  G�      F      ��  u vdd       F      �d  u vdd       F        u vdd       F        B�        �j  (� vdd       F        B�        �  (� vdd       F        B�        �  (� vdd       F        B�        �D  (� vdd       F        B�        �  (� vdd       F        B�        
�  (� vdd       F      �  u vdd       F      �(  u vdd       F      ��  z] 
vctrp       G   , �  d� �  f:   f:   d� �  d�      G   , ��  �� ��  �� ��  �� ��  �� ��  ��      G   , �  �� �  �x �  �x �  �� �  ��      G   , 	  �� 	  �x �  �x �  �� 	  ��      G   , �/  �� �/  ��    ��    �� �/  ��      G   , �.  �� �.  �x �  �x �  �� �.  ��      G   , k  �� k  �� S  �� S  �� k  ��      G   , �U  �� �U  �x �=  �x �=  �� �U  ��      G   , ��  �� ��  �x �y  �x �y  �� ��  ��      G   , ��  �� ��  �� ��  �� ��  �� ��  ��      G   ,  �  ��  �  �x  p  �x  p  ��  �  ��      G   ,  �  ��  �  ��  �  ��  �  ��  �  ��      G   , �a  S\ �a  V| �=  V| �=  S\ �a  S\      G   , #�  K� #�  M 'Y  M 'Y  K� #�  K�      G   , #�  P� #�  RD 'Y  RD 'Y  P� #�  P�   	   G   !     � $ F  f: F  � L  � L  �   	   G   !     �  _  �� _   &   	   G   !     �  �  �� �   &   	   G   !     �  �#  �� �#   &   	   G   !     �  ��  �� ��   &   	   G   !     �  ��  �� ��   &   	   G   !     �  �I  �� �I   &   	   G   !     �  ��  �� ��   &   	   G   !     �  �"  �� �"   &   	   G   !     � $ R�  � R�  # %�  # %�  R0   	   G   !     ,  � m� � R� �k R�   	   G   !     �  �O R� �O  T�   	   G   !     �  p� \d  � \d   	   G   !     ,  p\ m� p\ Zp   	   G   !     ,  e� m� e� Zp   	   G   !     ,  Z� m� Z� Zp   	   G   !     ,  P m� P Zp   	   G   !     ,  E< m� E< Zp   	   G   !     ,  :t m� :t Zp   	   G   !     ,  /� m� /� Zp   	   G   !     ,  $� m� $� Zp   	   G   !     ,   m�  Zp   	   G   !     ,  T m� T Zp   	   G   !     ,  � m� � Zp   	   G   !     ,   �� m�  �� Zp   	   G   !     ,   �� m�  �� Zp   	   G   !     ,   �4 m�  �4 Zp   	   G   !     ,   �l m�  �l Zp   	   G   !     ,   Τ m�  Τ Zp   	   G   !     ,   �� m�  �� Zp   	   G   !     ,   � m�  � Zp   	   G   !     ,   �L m�  �L Zp   	   G   !     ,   �� m�  �� Zp   	   G   !     ,   �� m�  �� Zp   	   G   !     ,   �� m�  �� Zp   	   G   !     ,   �, m�  �, Zp   	   G   !     ,   xd m�  xd Zp   	   G   !     �  �  �� �   &      G   , �  N* �  O� �  O� �  N* �  N*      G   , ��  N* ��  O� �y  O� �y  N* ��  N*      G   , �U  N* �U  O� �=  O� �=  N* �U  N*      G   , k  |. k  �� S  �� S  |. k  |.      G   , k  |. k  �� S  �� S  |. k  |.      G   , �/  |. �/  ��    ��    |. �/  |.      G   , �/  |. �/  ��    ��    |. �/  |.      G   , ��  |. ��  �� ��  �� ��  |. ��  |.      G   , ��  |. ��  �� ��  �� ��  |. ��  |.      G   , ��  |. ��  �� ��  �� ��  |. ��  |.      G   , ��  |. ��  �� ��  �� ��  |. ��  |.      G   , ��   & ��  !� ��  !� ��   & ��   &      G   , ��   & ��  !� ��  !� ��   & ��   &      G   , ��   & ��  !� ��  !� ��   & ��   &      G   , ��   & ��  !� ��  !� ��   & ��   &      G   , k   & k  !� S  !� S   & k   &      G   , k   & k  !� S  !� S   & k   &      G   , �/   & �/  !�    !�     & �/   &      G   , �/   & �/  !�    !�     & �/   &      G   , k  p! k  qk S  qk S  p! k  p!      G   ,   W   X\ �  X\ �  W   W      G   , ��  S� ��  U� �y  U� �y  S� ��  S�      G   , ��  G� ��  I� �y  I� �y  G� ��  G�      G   , k  t k  v S  v S  t k  t      G   , �/  t �/  v    v    t �/  t      G   , �  S� �  U� �  U� �  S� �  S�      G   , ��  t ��  v ��  v ��  t ��  t      G   , �U  S� �U  U� �=  U� �=  S� �U  S�      G   , ��  '� ��  )� ��  )� ��  '� ��  '�      G   , ��  '� ��  )� ��  )� ��  '� ��  '�      G   , �U  G� �U  I� �=  I� �=  G� �U  G�      G   , k  '� k  )� S  )� S  '� k  '�      G   , �  G� �  I� �  I� �  G� �  G�      G   , �/  '� �/  )�    )�    '� �/  '�      G   ,  w� m�  w� q�  x� q�  x� m�  w� m�      G   ,  �� m�  �� q�  �� q�  �� m�  �� m�      G   ,  �^ m�  �^ q�  �� q�  �� m�  �^ m�      G   ,  �& m�  �& q�  �R q�  �R m�  �& m�      G   ,  �� m�  �� q�  � q�  � m�  �� m�      G   ,  �� m�  �� q�  �� q�  �� m�  �� m�      G   ,  �~ m�  �~ q�  �� q�  �� m�  �~ m�      G   ,  �F m�  �F q�  �r q�  �r m�  �F m�      G   ,  � m�  � q�  �: q�  �: m�  � m�      G   ,  �� m�  �� q�  � q�  � m�  �� m�      G   ,  � m�  � q�  �� q�  �� m�  � m�      G   ,  �f m�  �f q�  � q�  � m�  �f m�      G   ,  �. m�  �. q�  �Z q�  �Z m�  �. m�      G   , � m� � q� " q� " m� � m�      G   , � m� � q� � q� � m� � m�      G   , � m� � q� � q� � m� � m�      G   , $N m� $N q� %z q� %z m� $N m�      G   , / m� / q� 0B q� 0B m� / m�      G   , 9� m� 9� q� ;
 q� ;
 m� 9� m�      G   , D� m� D� q� E� q� E� m� D� m�      G   , On m� On q� P� q� P� m� On m�      G   , Z6 m� Z6 q� [b q� [b m� Z6 m�      G   , d� m� d� q� f* q� f* m� d� m�      G   , o� m� o� q� p� q� p� m� o� m�      G   , z� m� z� q� {� q� {� m� z� m�      G   , �V m� �V q� �� q� �� m� �V m�      G   , � m� � q� �J q� �J m� � m�      G   , �� m� �� q� � q� � m� �� m�      G   , �� m� �� q� �� q� �� m� �� m�      G   , �v m� �v q� �� q� �� m� �v m�      G   , �> m� �> q� �j q� �j m� �> m�      G   , � m� � q� �2 q� �2 m� � m�      G   , �� m� �� q� �� q� �� m� �� m�      G   , ۖ m� ۖ q� �� q� �� m� ۖ m�      G   , �^ m� �^ q� � q� � m� �^ m�      G   , �& m� �& q� �R q� �R m� �& m�      G   , �� m� �� q� � q� � m� �� m�      G   , � m� � q� � q� � m� � m�      G   , ~ m� ~ q� � q� � m� ~ m�      G   , F m� F q� r q� r m� F m�      G   , ' m� ' q� (: q� (: m� ' m�      G   , 1� m� 1� q� 3 q� 3 m� 1� m�      G   , <� m� <� q� =� q� =� m� <� m�      G   ,  �  �  � ^X  � ^X  �  �  �  �      G   ,  �  �  � ^X  p ^X  p  �  �  �      G   ,  @�      @�  �  D>  �  D>      @�          G   ,  �2      �2  �  ��  �  ��      �2          G   ,  ת      ת  �  �.  �  �.      ת          G   , #"     #"  � &�  � &�     #"          G   , n�     n�  � r  � r     n�          G   , �     �  � ��  � ��     �          G   , �     �  � 	  � 	     �          G   , Q     Q  � T�  � T�     Q          F  , , �K  �; �K  � �  � �  �; �K  �;      F  , , �K  �� �K  �� �  �� �  �� �K  ��      F  , , �K  �[ �K  �# �  �# �  �[ �K  �[      F  , , �K  �� �K  �� �  �� �  �� �K  ��      F  , , �K  �{ �K  �C �  �C �  �{ �K  �{      F  , , �  �; �  � �  � �  �; �  �;      F  , , �  �� �  �� �  �� �  �� �  ��      F  , , �  �[ �  �# �  �# �  �[ �  �[      F  , , �  �� �  �� �  �� �  �� �  ��      F  , , �  �{ �  �C �  �C �  �{ �  �{      F  , , %  � %  �� �  �� �  � %  �      F  , , %  �� %  �d �  �d �  �� %  ��      F  , , %  �, %  �� �  �� �  �, %  �,      F  , , %  �� %  �� �  �� �  �� %  ��      F  , , %  �L %  � �  � �  �L %  �L      F  , , �  � �  �� ]  �� ]  � �  �      F  , , �  �� �  �d ]  �d ]  �� �  ��      F  , , �  �, �  �� ]  �� ]  �, �  �,      F  , , �  �� �  �� ]  �� ]  �� �  ��      F  , , �  �L �  � ]  � ]  �L �  �L      F  , , a  � a  �� )  �� )  � a  �      F  , , a  �� a  �d )  �d )  �� a  ��      F  , , a  �, a  �� )  �� )  �, a  �,      F  , , a  �� a  �� )  �� )  �� a  ��      F  , , a  �L a  � )  � )  �L a  �L      F  , , �  � �  �� �  �� �  � �  �      F  , , �  �� �  �d �  �d �  �� �  ��      F  , , �  �, �  �� �  �� �  �, �  �,      F  , , �  �� �  �� �  �� �  �� �  ��      F  , , �  �L �  � �  � �  �L �  �L      F  , , ��  �; ��  � �O  � �O  �; ��  �;      F  , , ��  �� ��  �� �O  �� �O  �� ��  ��      F  , , ��  �[ ��  �# �O  �# �O  �[ ��  �[      F  , , ��  �� ��  �� �O  �� �O  �� ��  ��      F  , , ��  �{ ��  �C �O  �C �O  �{ ��  �{      F  , , ��  �; ��  � ��  � ��  �; ��  �;      F  , , ��  �� ��  �� ��  �� ��  �� ��  ��      F  , , ��  �[ ��  �# ��  �# ��  �[ ��  �[      F  , , ��  �� ��  �� ��  �� ��  �� ��  ��      F  , , ��  �{ ��  �C ��  �C ��  �{ ��  �{      F  , , ׆  � ׆  �� �N  �� �N  � ׆  �      F  , , ׆  �� ׆  �d �N  �d �N  �� ׆  ��      F  , , ׆  �, ׆  �� �N  �� �N  �, ׆  �,      F  , , ׆  �� ׆  �� �N  �� �N  �� ׆  ��      F  , , ׆  �L ׆  � �N  � �N  �L ׆  �L      F  , , ��  � ��  �� ־  �� ־  � ��  �      F  , , ��  �� ��  �d ־  �d ־  �� ��  ��      F  , , ��  �, ��  �� ־  �� ־  �, ��  �,      F  , , ��  �� ��  �� ־  �� ־  �� ��  ��      F  , , ��  �L ��  � ־  � ־  �L ��  �L      F  , , �  �; �  � �  � �  �; �  �;      F  , , �  �� �  �� �  �� �  �� �  ��      F  , , �  �[ �  �# �  �# �  �[ �  �[      F  , , �  �� �  �� �  �� �  �� �  ��      F  , , �  �{ �  �C �  �C �  �{ �  �{      F  , , 3  �; 3  � �  � �  �; 3  �;      F  , , 3  �� 3  �� �  �� �  �� 3  ��      F  , , 3  �[ 3  �# �  �# �  �[ 3  �[      F  , , 3  �� 3  �� �  �� �  �� 3  ��      F  , , 3  �{ 3  �C �  �C �  �{ 3  �{      F  , , �  � �  �� �u  �� �u  � �  �      F  , , �  �� �  �d �u  �d �u  �� �  ��      F  , , �  �, �  �� �u  �� �u  �, �  �,      F  , , �  �� �  �� �u  �� �u  �� �  ��      F  , , �  �L �  � �u  � �u  �L �  �L      F  , , �  � �  �� ��  �� ��  � �  �      F  , , �  �� �  �d ��  �d ��  �� �  ��      F  , , �  �, �  �� ��  �� ��  �, �  �,      F  , , �  �� �  �� ��  �� ��  �� �  ��      F  , , �  �L �  � ��  � ��  �L �  �L      F  , , ��  � ��  �� ��  �� ��  � ��  �      F  , , ��  �� ��  �d ��  �d ��  �� ��  ��      F  , , ��  �, ��  �� ��  �� ��  �, ��  �,      F  , , ��  �� ��  �� ��  �� ��  �� ��  ��      F  , , ��  �L ��  � ��  � ��  �L ��  �L      F  , , �Y  � �Y  �� �!  �� �!  � �Y  �      F  , , �Y  �� �Y  �d �!  �d �!  �� �Y  ��      F  , , �Y  �, �Y  �� �!  �� �!  �, �Y  �,      F  , , �Y  �� �Y  �� �!  �� �!  �� �Y  ��      F  , , �Y  �L �Y  � �!  � �!  �L �Y  �L      F  , , �3  �; �3  � ��  � ��  �; �3  �;      F  , , �3  �� �3  �� ��  �� ��  �� �3  ��      F  , , �3  �[ �3  �# ��  �# ��  �[ �3  �[      F  , , �3  �� �3  �� ��  �� ��  �� �3  ��      F  , , �3  �{ �3  �C ��  �C ��  �{ �3  �{      F  , , ݣ  �; ݣ  � �k  � �k  �; ݣ  �;      F  , , ݣ  �� ݣ  �� �k  �� �k  �� ݣ  ��      F  , , ݣ  �[ ݣ  �# �k  �# �k  �[ ݣ  �[      F  , , ݣ  �� ݣ  �� �k  �� �k  �� ݣ  ��      F  , , ݣ  �{ ݣ  �C �k  �C �k  �{ ݣ  �{      F  , , �  e �  e� r  e� r  e �  e      F  , ,   e   e� �  e� �  e   e      F  , , �{  S� �{  T� �C  T� �C  S� �{  S�      F  , , �{  UP �{  V �C  V �C  UP �{  UP      F  , , ��  S� ��  T� ȳ  T� ȳ  S� ��  S�      F  , , ��  UP ��  V ȳ  V ȳ  UP ��  UP      F  , , �[  S� �[  T� �#  T� �#  S� �[  S�      F  , , �[  UP �[  V �#  V �#  UP �[  UP      F  , , %�  K� %�  L� &�  L� &�  K� %�  K�      F  , , $k  K� $k  L� %3  L� %3  K� $k  K�      F  , , %�  Q" %�  Q� &�  Q� &�  Q" %�  Q"      F  , , $k  Q" $k  Q� %3  Q� %3  Q" $k  Q"      F  , ,  $  �  $  ��  �  ��  �  �  $  �      F  , ,  $  ��  $  �d  �  �d  �  ��  $  ��      F  , ,  $  �,  $  ��  �  ��  �  �,  $  �,      F  , ,  $  ��  $  ��  �  ��  �  ��  $  ��      F  , ,  $  �L  $  �  �  �  �  �L  $  �L      F  , ,  �  �  �  ��  \  ��  \  �  �  �      F  , ,  �  ��  �  �d  \  �d  \  ��  �  ��      F  , ,  �  �,  �  ��  \  ��  \  �,  �  �,      F  , ,  �  ��  �  ��  \  ��  \  ��  �  ��      F  , ,  �  �L  �  �  \  �  \  �L  �  �L      F  , ,    �    ��  �  ��  �  �    �      F  , ,    ��    �d  �  �d  �  ��    ��      F  , ,    �,    ��  �  ��  �  �,    �,      F  , ,    ��    ��  �  ��  �  ��    ��      F  , ,    �L    �  �  �  �  �L    �L      F  , ,  
�  �;  
�  �  T  �  T  �;  
�  �;      F  , ,  
�  ��  
�  ��  T  ��  T  ��  
�  ��      F  , ,  
�  �[  
�  �#  T  �#  T  �[  
�  �[      F  , ,  
�  ��  
�  ��  T  ��  T  ��  
�  ��      F  , ,  
�  �{  
�  �C  T  �C  T  �{  
�  �{      F  , ,  �  �;  �  �  	�  �  	�  �;  �  �;      F  , ,  �  ��  �  ��  	�  ��  	�  ��  �  ��      F  , ,  �  �[  �  �#  	�  �#  	�  �[  �  �[      F  , ,  �  ��  �  ��  	�  ��  	�  ��  �  ��      F  , ,  �  �{  �  �C  	�  �C  	�  �{  �  �{      F  , ,  l  �;  l  �  4  �  4  �;  l  �;      F  , ,  l  ��  l  ��  4  ��  4  ��  l  ��      F  , ,  l  �[  l  �#  4  �#  4  �[  l  �[      F  , ,  l  ��  l  ��  4  ��  4  ��  l  ��      F  , ,  l  �{  l  �C  4  �C  4  �{  l  �{      F  , ,  �  �;  �  �  �  �  �  �;  �  �;      F  , ,  �  ��  �  ��  �  ��  �  ��  �  ��      F  , ,  �  �[  �  �#  �  �#  �  �[  �  �[      F  , ,  �  ��  �  ��  �  ��  �  ��  �  ��      F  , ,  �  �{  �  �C  �  �C  �  �{  �  �{      F  , ,  L  �;  L  �    �    �;  L  �;      F  , ,  L  ��  L  ��    ��    ��  L  ��      F  , ,  L  �[  L  �#    �#    �[  L  �[      F  , ,  L  ��  L  ��    ��    ��  L  ��      F  , ,  L  �{  L  �C    �C    �{  L  �{      F  , ,  D  �  D  ��    ��    �  D  �      F  , ,  D  ��  D  �d    �d    ��  D  ��      F  , ,  D  �,  D  ��    ��    �,  D  �,      F  , ,  D  ��  D  ��    ��    ��  D  ��      F  , ,  D  �L  D  �    �    �L  D  �L      F  , ,  �  �  �  ��  |  ��  |  �  �  �      F  , ,  �  ��  �  �d  |  �d  |  ��  �  ��      F  , ,  �  �,  �  ��  |  ��  |  �,  �  �,      F  , ,  �  ��  �  ��  |  ��  |  ��  �  ��      F  , ,  �  �L  �  �  |  �  |  �L  �  �L      F  , , �Y  T� �Y  UP �!  UP �!  T� �Y  T�      F  , , �Y  H� �Y  I\ �!  I\ �!  H� �Y  H�      F  , , 3  t� 3  ul �  ul �  t� 3  t�      F  , , ��  t� ��  ul ��  ul ��  t� ��  t�      F  , , �  T� �  UP ]  UP ]  T� �  T�      F  , , �  t� �  ul �  ul �  t� �  t�      F  , , �  T� �  UP ��  UP ��  T� �  T�      F  , , �  (x �  )@ �  )@ �  (x �  (x      F  , , ݣ  (x ݣ  )@ �k  )@ �k  (x ݣ  (x      F  , , �  H� �  I\ ��  I\ ��  H� �  H�      F  , , 3  (x 3  )@ �  )@ �  (x 3  (x      F  , , �  H� �  I\ ]  I\ ]  H� �  H�      F  , , ��  (x ��  )@ ��  )@ ��  (x ��  (x      F  , , ��  T� ��  UP ��  UP ��  T� ��  T�      F  , , ��  H� ��  I\ ��  I\ ��  H� ��  H�      F  , , �  t� �  ul �  ul �  t� �  t�      F  , , ��  t� ��  ul �O  ul �O  t� ��  t�      F  , , %  T� %  UP �  UP �  T� %  T�      F  , , �K  t� �K  ul �  ul �  t� �K  t�      F  , , �  T� �  UP �u  UP �u  T� �  T�      F  , , �K  (x �K  )@ �  )@ �  (x �K  (x      F  , , �3  (x �3  )@ ��  )@ ��  (x �3  (x      F  , , �  H� �  I\ �u  I\ �u  H� �  H�      F  , , �  (x �  )@ �  )@ �  (x �  (x      F  , , %  H� %  I\ �  I\ �  H� %  H�      F  , , ��  (x ��  )@ �O  )@ �O  (x ��  (x      F  , , 3  pb 3  q* �  q* �  pb 3  pb      F  , , �  pb �  q* �  q* �  pb �  pb      F  , , �  N� �  OV ]  OV ]  N� �  N�      F  , , �Y  N� �Y  OV �!  OV �!  N� �Y  N�      F  , , �  N� �  OV ��  OV ��  N� �  N�      F  , , 3  |� 3  }Z �  }Z �  |� 3  |�      F  , , 3  |� 3  }Z �  }Z �  |� 3  |�      F  , , ��  |� ��  }Z ��  }Z ��  |� ��  |�      F  , , ��  |� ��  }Z ��  }Z ��  |� ��  |�      F  , , �  |� �  }Z �  }Z �  |� �  |�      F  , , �  |� �  }Z �  }Z �  |� �  |�      F  , , ݣ  |� ݣ  }Z �k  }Z �k  |� ݣ  |�      F  , , ݣ  |� ݣ  }Z �k  }Z �k  |� ݣ  |�      F  , , �   � �  !R �  !R �   � �   �      F  , , �   � �  !R �  !R �   � �   �      F  , , ݣ   � ݣ  !R �k  !R �k   � ݣ   �      F  , , ݣ   � ݣ  !R �k  !R �k   � ݣ   �      F  , , 3   � 3  !R �  !R �   � 3   �      F  , , 3   � 3  !R �  !R �   � 3   �      F  , , ��   � ��  !R ��  !R ��   � ��   �      F  , , ��   � ��  !R ��  !R ��   � ��   �      F  , , %  N� %  OV �  OV �  N� %  N�      F  , , ��  N� ��  OV ��  OV ��  N� ��  N�      F  , , �  N� �  OV �u  OV �u  N� �  N�      F  , , �  |� �  }Z �  }Z �  |� �  |�      F  , , �  |� �  }Z �  }Z �  |� �  |�      F  , , ��  |� ��  }Z �O  }Z �O  |� ��  |�      F  , , ��  |� ��  }Z �O  }Z �O  |� ��  |�      F  , , �K  |� �K  }Z �  }Z �  |� �K  |�      F  , , �K  |� �K  }Z �  }Z �  |� �K  |�      F  , , �3  |� �3  }Z ��  }Z ��  |� �3  |�      F  , , �3  |� �3  }Z ��  }Z ��  |� �3  |�      F  , , �K   � �K  !R �  !R �   � �K   �      F  , , �K   � �K  !R �  !R �   � �K   �      F  , , �3   � �3  !R ��  !R ��   � �3   �      F  , , �3   � �3  !R ��  !R ��   � �3   �      F  , , �   � �  !R �  !R �   � �   �      F  , , �   � �  !R �  !R �   � �   �      F  , , ��   � ��  !R �O  !R �O   � ��   �      F  , , ��   � ��  !R �O  !R �O   � ��   �      F  , , �  WS �  X �  X �  WS �  WS      F  , , �  WS �  X T  X T  WS �  WS      D   , �  d� �  f:   f:   d� �  d�   	   D   !       �N  ^� �  ^�   	   D   !       և  >� �  >�   	   D   !     �  �F  |� �  |�   	   D   !     �  �z  N� �F  N� �F  N�   	   D   !     �  �)   � �   �   	   D   !     �  �T  |� �  |�   	   D   !     �  �   � �T   �   	   D   !     r  �q  Q� �q  N*   	   D   !     r  �  Q� �  N*   	   D   !     r   �  Q�  �  N*   	   D   !     r  �  K� �  O�   	   D   !     r  �]  K� �]  O�   	   D   !     r  ��  K� ��  O�   	   D   !     r  ��  K� ��  O�   	   D   !     r  7  K� 7  O�   	   D   !     r  
�  K� 
�  O�   	   D   !     r  K  Q� K  N*   	   D   !     r  ��  Q� ��  N*   	   D   !     r  �]  Q� �]  N*   	   D   !     r  ��  Q� ��  N*   	   D   !     r  ��  Q� ��  N*   	   D   !     r  ��  K� ��  O�   	   D   !     r  �q  K� �q  O�   	   D   !     r  �  K� �  O�   	   D   !     r   �  K�  �  O�   	   D   !     r  K  K� K  O�   	   D   !     r  �  K� �  O�   	   D   !     r  7  Q� 7  N*   	   D   !     r  �  Q� �  N*   	   D   !     �  �  N� �  N�   	   D   !     �  �T  N� �  N�   	   D   !     �  �  N� �T  N�   	   D   !     �  �z  N� �  N�   	   D   !     �  �  N� �  N�   	   D   !     �  �  N� �T  N�   	   D   !     �  �T  N� �  N�   	   D   !     �  �  N� 	�  N�   	   D   !     �  	�  N� .  N�   	   D   !     �  	�  N� �  N�   	   D   !     �  �  N� �z  N�   	   D   !     @  �T  b �W  b   	   D   !     @  ��  ;� �T  ;�   	   D   !     �  	�  |� �  |�   	   D   !      �  ��  \� ��  S�   	   D   !      �  |  \� |  S�   	   D   !      �  �  o a  o   	   D   !     �  �  |� �T  |�   	   D   !     @  �  b ��  b   	   D   !     @  	�  b �  b   	   D   !     @  ��  b �T  b   	   D   !     @  �  b �  b   	   D   !     r   �  }�  �  y�   	   D   !     r  K  }� K  y�   	   D   !     r  ��  }� ��  y�   	   D   !     r  7  }� 7  y�   	   D   !      �  ��  xi ��  f�   	   D   !      �  |  xi |  f�   	   D   !     @  	�  b   b �  b   	   D   !       �  e� �  e�   	   D   !       �  e� 	  e�   	   D   !      �  �@  \� �@  S�   	   D   !     r  �]  }� �]  y�   	   D   !     r  ��  }� ��  y�   	   D   !      �  �  \� �  S�   	   D   !     @  �  b �  b   	   D   !     @  �z  b �/  b   	   D   !     r  �  }� �  y�   	   D   !      �  �  xi �  f�   	   D   !      �  �@  xi �@  f�   	   D   !     @  �  b �z  b   	   D   !     r  �q  }� �q  y�   	   D   !      �  �  xi �  f�   	   D   !     �  �  |� �  |�   	   D   !     @  �  b �  b   	   D   !     @  �  b �  b   	   D   !     @  �J  b �  b   	   D   !     r  ��  }� ��  y�   	   D   !     �  �  |� �z  |�   	   D   !     r  �  }� �  y�   	   D   !      �  �  \� �  S�   	   D   !     @  �  ;� �  ;�   	   D   !     @  �  ;� ��  ;�   	   D   !     @  �z  ;� �/  ;�   	   D   !     r  ��   & ��  #�   	   D   !     �  �z   � �   �   	   D   !     �  �   � �   �   	   D   !     r  �q   & �q  #�   	   D   !     @  �  ;� �  ;�   	   D   !     r  �   & �  #�   	   D   !     r  �]   & �]  #�   	   D   !     r  ��   & ��  #�   	   D   !     @  �"  ;� �  ;�   	   D   !      �  �  @� �  J=   	   D   !      �  �,  @� �,  J=   	   D   !      �  �  %{ �  6�   	   D   !      �  ��  @� ��  J=   	   D   !      �  ��  %{ ��  6�   	   D   !      �  �,  %{ �,  6�   	   D   !     r  �   & �  #�   	   D   !     @  �z  ;� �w  ;�   	   D   !     �  	�   � .   �   	   D   !     @  �  ;� .  ;�   	   D   !     r  ��   & ��  #�   	   D   !     r  7   & 7  #�   	   D   !     r  
�   & 
�  #�   	   D   !     @  	�  ;� �  ;�   	   D   !     @  �  ;� .  ;�   	   D   !     @  �T  ;� �Q  ;�   	   D   !     r   �   &  �  #�   	   D   !      �  �h  @� �h  J=   	   D   !      �    @�   J=   	   D   !      �  �  @� �  J=   	   D   !     r  K   & K  #�   	   D   !      �  �h  %{ �h  6�   	   D   !      �    %{   6�   	   D   !      �  �  %{ �  6�   	   D   !     @  �  ;� �  ;�   	   D   !     r  �   & �  #�   	   D   !     @  �^  ;� �  ;�   	   D   !     @  �  ;� 	�  ;�   	   D   !     �  �T   � �   �   	   D   !     �  �   � 	�   �      D   , ��  N* ��  O� �z  O� �z  N* ��  N*      D   , �F  N* �F  O� ��  O� ��  N* �F  N*      D   , �  N* �  O� �  O� �  N* �  N*      D   , ��  N* ��  O� �y  O� �y  N* ��  N*      D   , �U  N* �U  O� �=  O� �=  N* �U  N*      D   , �  |. �  }� �T  }� �T  |. �  |.      D   , �   & �  !� �T  !� �T   & �   &      D   , �  N* �  O� �  O� �  N* �  N*      D   , �  N* �  O� �T  O� �T  N* �  N*      D   , �T  N* �T  O� �  O� �  N* �T  N*      D   , �z  N* �z  O� �  O� �  N* �z  N*      D   , �  N* �  O� �  O� �  N* �  N*      D   , �  N* �  O� �T  O� �T  N* �  N*      D   , �T  N* �T  O� �  O� �  N* �T  N*      D   , �  N* �  O� 	�  O� 	�  N* �  N*      D   , 	�  N* 	�  O� .  O� .  N* 	�  N*      D   , �  N* �  O� 	�  O� 	�  N* �  N*      D   , �z  N* �z  O� �  O� �  N* �z  N*      D   , ��  y� ��  { �>  { �>  y� ��  y�      D   , ��  y� ��  z� �>  z� �>  y� ��  y�      D   , ��  P� ��  R0 �>  R0 �>  P� ��  P�      D   , ��  Q ��  Q� �>  Q� �>  Q ��  Q      D   , ��  K� ��  L� �>  L� �>  K� ��  K�      D   , ��  K� ��  L� �>  L� �>  K� ��  K�      D   , ��  "� ��  $, �>  $, �>  "� ��  "�      D   , ��  # ��  #� �>  #� �>  # ��  #      D   , �  |. �  }� 	�  }� 	�  |. �  |.      D   ,   y�   { z  { z  y�   y�      D   ,   y�   z� z  z� z  y�   y�      D   ,   Q   Q� z  Q� z  Q   Q      D   ,   P�   R0 z  R0 z  P�   P�      D   , f  f� f  m� �  m� �  f� f  f�      D   , M  t M  v �  v �  t M  t      D   , �  t �  v 
I  v 
I  t �  t      D   , �  y� �  z� 	  z� 	  y� �  y�      D   , %  n� %  o� e  o� e  n� %  n�      D   , *  g *  h j  h j  g *  g      D   , �  l� �  m� ,  m� ,  l� �  l�      D   , p  l� p  m� �  m� �  l� p  l�      D   , �  f� �  g� �  g� �  f� �  f�      D   , 2  f� 2  g� r  g� r  f� 2  f�      D   , -  f� -  g� w  g� w  f� -  f�      D   , �  f� �  g� �  g� �  f� �  f�      D   , �  n} �  o� �  o� �  n} �  n}      D   , �  f� �  m� �  m� �  f� �  f�      D   , _  f� _  m� E  m� E  f� _  f�      D   , �  f� �  m� �  m� �  f� �  f�      D   ,   f�   m� �  m� �  f�   f�      D   ,   f�   m� �  m� �  f�   f�      D   , �  f� �  m� �  m� �  f� �  f�      D   , �  f� �  m� �  m� �  f� �  f�      D   , W  f� W  m� =  m� =  f� W  f�      D   , 	  q� 	  xi 
  xi 
  q� 	  q�      D   , �  p5 �  qW �  qW �  p5 �  p5      D   , �  q� �  xi y  xi y  q� �  q�      D   , �  q� �  xi y  xi y  q� �  q�      D   , �  f� �  m� y  m� y  f� �  f�      D   , #  p? #  qM ~  qM ~  p? #  p?      D   , k  |. k  }� S  }� S  |. k  |.      D   , k  |. k  }� S  }� S  |. k  |.      D   , ��  t ��  v �  v �  t ��  t      D   , �k  q� �k  xi �Q  xi �Q  q� �k  q�      D   , 	  q� 	  xi �  xi �  q� 	  q�      D   , �j  y� �j  z� ��  z� ��  y� �j  y�      D   , ��  t ��  v �  v �  t ��  t      D   , �j  y� �j  { ��  { ��  y� �j  y�      D   ,   q�   xi e  xi e  q�   q�      D   , �T  |. �T  }� �  }� �  |. �T  |.      D   , ��  q� ��  xi ��  xi ��  q� ��  q�      D   , �k  q� �k  xi �Q  xi �Q  q� �k  q�      D   , ��  y� ��  z� f  z� f  y� ��  y�      D   , 	  q� 	  xi �  xi �  q� 	  q�      D   , ��  f� ��  m� ��  m� ��  f� ��  f�      D   ,   q�   xi e  xi e  q�   q�      D   , �k  f� �k  m� �Q  m� �Q  f� �k  f�      D   , 	  f� 	  m� �  m� �  f� 	  f�      D   , 9  t 9  v �  v �  t 9  t      D   , ��  y� ��  z� �R  z� �R  y� ��  y�      D   , ��  f� ��  m�    m�    f� ��  f�      D   , 9  t 9  v �  v �  t 9  t      D   , ��  q� ��  xi ��  xi ��  q� ��  q�      D   , ��  q� ��  xi ��  xi ��  q� ��  q�      D   , �W  q� �W  xi �=  xi �=  q� �W  q�      D   , �V  y� �V  z� ��  z� ��  y� �V  y�      D   , �W  f� �W  m� �=  m� �=  f� �W  f�      D   , �  t �  v ��  v ��  t �  t      D   , �*  f� �*  m� �j  m� �j  f� �*  f�      D   , �W  q� �W  xi �=  xi �=  q� �W  q�      D   , ~  y� ~  z� �  z� �  y� ~  y�      D   , ��  q� ��  xi ��  xi ��  q� ��  q�      D   , ��  t ��  v  !  v  !  t ��  t      D   , �/  |. �/  }�    }�    |. �/  |.      D   , �/  |. �/  }�    }�    |. �/  |.      D   , R  Zs R  \� �  \� �  Zs R  Zs      D   ,   S�   V1 e  V1 e  S�   S�      D   , ��  Q ��  Q� f  Q� f  Q ��  Q      D   , ��  S� ��  U� �  U� �  S� ��  S�      D   , �k  S� �k  V1 �Q  V1 �Q  S� �k  S�      D   , ��  Zs ��  \� ��  \� ��  Zs ��  Zs      D   , ��  S� ��  V1 ��  V1 ��  S� ��  S�      D   , 	  S� 	  V1 �  V1 �  S� 	  S�      D   , ��  al ��  b�    b�    al ��  al      D   , ��  Zs ��  \�    \�    Zs ��  Zs      D   , 9  S� 9  U� �  U� �  S� 9  S�      D   , �k  Zs �k  \� �Q  \� �Q  Zs �k  Zs      D   , ��  Q ��  Q� �R  Q� �R  Q ��  Q      D   , 	  Zs 	  \� �  \� �  Zs 	  Zs      D   , ~  Q ~  Q� �  Q� �  Q ~  Q      D   , ��  al ��  b� ��  b� ��  al ��  al      D   , <  al <  b� �  b� �  al <  al      D   ,   S�   V1 e  V1 e  S�   S�      D   , ��  S� ��  V1 ��  V1 ��  S� ��  S�      D   , ��  S� ��  U�  !  U�  !  S� ��  S�      D   , �j  P� �j  R0 ��  R0 ��  P� �j  P�      D   , ��  S� ��  U� �  U� �  S� ��  S�      D   , ��  Zs ��  \� ��  \� ��  Zs ��  Zs      D   , ��  Zs ��  \� ��  \� ��  Zs ��  Zs      D   , ��  S� ��  V1 ��  V1 ��  S� ��  S�      D   , �k  S� �k  V1 �Q  V1 �Q  S� �k  S�      D   , 9  S� 9  U� �  U� �  S� 9  S�      D   , 	  S� 	  V1 �  V1 �  S� 	  S�      D   , �  S� �  U� ��  U� ��  S� �  S�      D   , �W  S� �W  V1 �=  V1 �=  S� �W  S�      D   , �W  Zs �W  \� �=  \� �=  Zs �W  Zs      D   , ��  ^t ��  _� \  _� \  ^t ��  ^t      D   , �*  al �*  b� �j  b� �j  al �*  al      D   , �*  Zs �*  \� �j  \� �j  Zs �*  Zs      D   , �V  Q �V  Q� ��  Q� ��  Q �V  Q      D   , �W  Zs �W  \� �=  \� �=  Zs �W  Zs      D   , �W  S� �W  V1 �=  V1 �=  S� �W  S�      D   , �j  Q �j  Q� ��  Q� ��  Q �j  Q      D   , ��  Zs ��  \� ��  \� ��  Zs ��  Zs      D   ,   Zs   \� e  \� e  Zs   Zs      D   , ��  S� ��  V1 ��  V1 ��  S� ��  S�      D   , �  S� �  U� 
I  U� 
I  S� �  S�      D   , �  Zs �  \� 
0  \� 
0  Zs �  Zs      D   , 	  S� 	  V1 
  V1 
  S� 	  S�      D   , �  a� �  b� 7  b� 7  a� �  a�      D   , �  e �  f �  f �  e �  e      D   , 2  e 2  f r  f r  e 2  e      D   , *  [� *  \� j  \� j  [� *  [�      D   , 2  [� 2  \� r  \� r  [� 2  [�      D   , -  d� -  f w  f w  d� -  d�      D   , 	  Zs 	  \� 
  \� 
  Zs 	  Zs      D   , �  Q �  Q� 	  Q� 	  Q �  Q      D   , �  Zs �  \� y  \� y  Zs �  Zs      D   , f  al f  b� �  b� �  al f  al      D   , �  Zs �  \� y  \� y  Zs �  Zs      D   ,   W0   X> y  X> y  W0   W0      D   , ]  al ]  b� �  b� �  al ]  al      D   , M  S� M  U� �  U� �  S� M  S�      D   , �  S� �  V1 y  V1 y  S� �  S�      D   , f  Zs f  \� �  \� �  Zs f  Zs      D   , �  S� �  V1 y  V1 y  S� �  S�      D   , �  d� �  f �  f �  d� �  d�      D   , �  [� �  \� �  \� �  [� �  [�      D   , �  Z� �  [� ,  [� ,  Z� �  Z�      D   , p  Z� p  [� �  [� �  Z� p  Z�      D   ,   Zs   \� �  \� �  Zs   Zs      D   , _  Zs _  \� E  \� E  Zs _  Zs      D   , �  W& �  XH �  XH �  W& �  W&      D   , �  Zs �  \� �  \� �  Zs �  Zs      D   , �  Zs �  \� �  \� �  Zs �  Zs      D   , W  Zs W  \� =  \� =  Zs W  Zs      D   , �  Zs �  \� �  \� �  Zs �  Zs      D   ,   Zs   \� �  \� �  Zs   Zs      D   , �  Zs �  \� �  \� �  Zs �  Zs      D   , �z  |. �z  }� �  }� �  |. �z  |.      D   , �  q� �  xi �w  xi �w  q� �  q�      D   , �  f� �  m� �w  m� �w  f� �  f�      D   , �  q� �  xi �w  xi �w  q� �  q�      D   , �  S� �  V1 �w  V1 �w  S� �  S�      D   , �  Zs �  \� �w  \� �w  Zs �  Zs      D   , �  S� �  V1 �w  V1 �w  S� �  S�      D   , �/  q� �/  xi �  xi �  q� �/  q�      D   , ��  q� ��  xi ��  xi ��  q� ��  q�      D   , �C  q� �C  xi �)  xi �)  q� �C  q�      D   , �B  y� �B  z� ��  z� ��  y� �B  y�      D   , �  q� �  xi �  xi �  q� �  q�      D   , �  q� �  xi �  xi �  q� �  q�      D   , �/  q� �/  xi �  xi �  q� �/  q�      D   , ��  q� ��  xi ��  xi ��  q� ��  q�      D   , �.  y� �.  z� �  z� �  y� �.  y�      D   , ��  f� ��  m� ��  m� ��  f� ��  f�      D   , �  q� �  xi �  xi �  q� �  q�      D   , �_  t �_  v ��  v ��  t �_  t      D   , �  f� �  m� ��  m� ��  f� �  f�      D   , �  q� �  xi �  xi �  q� �  q�      D   , �_  t �_  v ��  v ��  t �_  t      D   , ��  f� ��  m� �.  m� �.  f� ��  f�      D   , �  y� �  z� �  z� �  y� �  y�      D   , �  y� �  z� �  z� �  y� �  y�      D   , �  y� �  { �  { �  y� �  y�      D   , �  q� �  xi �  xi �  q� �  q�      D   , �  q� �  xi �  xi �  q� �  q�      D   , ��  t ��  v �o  v �o  t ��  t      D   , �  y� �  z� �  z� �  y� �  y�      D   , �.  y� �.  { �  { �  y� �.  y�      D   , ��  t ��  v �G  v �G  t ��  t      D   , �  f� �  m� �  m� �  f� �  f�      D   , ��  t ��  v �o  v �o  t ��  t      D   , �s  t �s  v ��  v ��  t �s  t      D   , �C  q� �C  xi �)  xi �)  q� �C  q�      D   , ��  |. ��  }� ��  }� ��  |. ��  |.      D   , ��  |. ��  }� ��  }� ��  |. ��  |.      D   , �  |. �  }� �  }� �  |. �  |.      D   , �  y� �  z� �*  z� �*  y� �  y�      D   , �  f� �  m� �  m� �  f� �  f�      D   , �/  f� �/  m� �  m� �  f� �/  f�      D   , ��  t ��  v �3  v �3  t ��  t      D   , �|  y� �|  z� ��  z� ��  y� �|  y�      D   , �  q� �  xi ��  xi ��  q� �  q�      D   , �F  |. �F  }� ��  }� ��  |. �F  |.      D   , ��  |. ��  }� �z  }� �z  |. ��  |.      D   , �P  y� �P  { ��  { ��  y� �P  y�      D   , �i  y� �i  { ��  { ��  y� �i  y�      D   , ��  |. ��  }� ��  }� ��  |. ��  |.      D   , ��  |. ��  }� ��  }� ��  |. ��  |.      D   , �}  q� �}  xi �c  xi �c  q� �}  q�      D   , �  q� �  xi ��  xi ��  q� �  q�      D   , �  y� �  z� �x  z� �x  y� �  y�      D   , �P  q� �P  xi �  xi �  q� �P  q�      D   , �  S� �  V1 ��  V1 ��  S� �  S�      D   , �(  P� �(  R0 �  R0 �  P� �(  P�      D   , �  P� �  R0 �s  R0 �s  P� �  P�      D   , ��  S� ��  U� �3  U� �3  S� ��  S�      D   , �5  S\ �5  T� ٧  T� ٧  S\ �5  S\      D   , �  Q �  Q� �x  Q� �x  Q �  Q      D   , ��  al ��  b� �  b� �  al ��  al      D   , �}  S� �}  V1 �c  V1 �c  S� �}  S�      D   , �  S� �  V1 ��  V1 ��  S� �  S�      D   , �N  ^t �N  _� َ  _� َ  ^t �N  ^t      D   , �P  S� �P  V1 �  V1 �  S� �P  S�      D   , �/  al �/  b� �o  b� �o  al �/  al      D   , �<  P� �<  R0 �  R0 �  P� �<  P�      D   , �  S� �  V1 �  V1 �  S� �  S�      D   , �  S� �  V1 �  V1 �  S� �  S�      D   , �  Q �  Q� �  Q� �  Q �  Q      D   , ��  Zs ��  \� �.  \� �.  Zs ��  Zs      D   , ��  S� ��  U� �G  U� �G  S� ��  S�      D   , �  Q �  Q� �  Q� �  Q �  Q      D   , �_  S� �_  U� ��  U� ��  S� �_  S�      D   , �_  S� �_  U� ��  U� ��  S� �_  S�      D   , �  Zs �  \� �  \� �  Zs �  Zs      D   , �/  S� �/  V1 �  V1 �  S� �/  S�      D   , �  Zs �  \� �  \� �  Zs �  Zs      D   , �  Zs �  \� �  \� �  Zs �  Zs      D   , �.  P� �.  R0 �  R0 �  P� �.  P�      D   , �.  P� �.  R0 �  R0 �  P� �.  P�      D   , �C  Zs �C  \� �)  \� �)  Zs �C  Zs      D   , ��  S� ��  U� �o  U� �o  S� ��  S�      D   , �  P� �  R0 �  R0 �  P� �  P�      D   , �/  S� �/  V1 �  V1 �  S� �/  S�      D   , ��  S� ��  V1 ��  V1 ��  S� ��  S�      D   , �  al �  b� ��  b� ��  al �  al      D   , �C  S� �C  V1 �)  V1 �)  S� �C  S�      D   , �  Zs �  \� �V  \� �V  Zs �  Zs      D   , �.  Q �.  Q� �  Q� �  Q �.  Q      D   , �  Q �  Q� �*  Q� �*  Q �  Q      D   , ��  S� ��  V1 ��  V1 ��  S� ��  S�      D   , �   al �   b� �J  b� �J  al �   al      D   , �C  S� �C  V1 �)  V1 �)  S� �C  S�      D   , �/  Zs �/  \� �  \� �  Zs �/  Zs      D   , �  Zs �  \� ��  \� ��  Zs �  Zs      D   , ��  Zs ��  \� ��  \� ��  Zs ��  Zs      D   , �  Zs �  \� �  \� �  Zs �  Zs      D   , �  S� �  V1 �  V1 �  S� �  S�      D   , �  P� �  R0 �  R0 �  P� �  P�      D   , ��  S� ��  U� �o  U� �o  S� ��  S�      D   , �  Q �  Q� �  Q� �  Q �  Q      D   , �b  al �b  b� �  b� �  al �b  al      D   , �B  Q �B  Q� ��  Q� ��  Q �B  Q      D   , ��  ^t ��  _� �   _� �   ^t ��  ^t      D   , �  S� �  V1 �  V1 �  S� �  S�      D   , �  S� �  V1 �  V1 �  S� �  S�      D   , �s  S� �s  U� ��  U� ��  S� �s  S�      D   , ��  al ��  b� �.  b� �.  al ��  al      D   , �x  Zs �x  \� �  \� �  Zs �x  Zs      D   , �  Zs �  \� �  \� �  Zs �  Zs      D   , �  S� �  V1 �  V1 �  S� �  S�      D   , �K  G� �K  I� �  I� �  G� �K  G�      D   , �d  ;8 �d  <x �  <x �  ;8 �d  ;8      D   , �  @� �  Cq �w  Cq �w  @� �  @�      D   , �  G� �  J= �w  J= �w  G� �  G�      D   , �  G� �  J= �w  J= �w  G� �  G�      D   , �d  @� �d  Cq �  Cq �  @� �d  @�      D   , �  @� �  Cq �w  Cq �w  @� �  @�      D   , �d  0/ �d  6� �  6� �  0/ �d  0/      D   , �  0/ �  6� �w  6� �w  0/ �  0/      D   , �z   & �z  !� �  !� �   & �z   &      D   , �  %{ �  ,= �w  ,= �w  %{ �  %{      D   , �  %{ �  ,= �w  ,= �w  %{ �  %{      D   , �K  '� �K  )� �  )� �  '� �K  '�      D   , ��  @� ��  Cq ��  Cq ��  @� ��  @�      D   , �  @� �  Cq �V  Cq �V  @� �  @�      D   , �  @� �  Cq �  Cq �  @� �  @�      D   , ��  G� ��  I� �o  I� �o  G� ��  G�      D   , �  K� �  L� �*  L� �*  K� �  K�      D   , �  G� �  J= �  J= �  G� �  G�      D   , �  G� �  J= �  J= �  G� �  G�      D   , ��  ;8 ��  <x ��  <x ��  ;8 ��  ;8      D   , �C  G� �C  J= �)  J= �)  G� �C  G�      D   , �.  K� �.  L� �  L� �  K� �.  K�      D   , �  >b �  ?p �  ?p �  >b �  >b      D   , �/  G� �/  J= �  J= �  G� �/  G�      D   , ��  @� ��  Cq ��  Cq ��  @� ��  @�      D   , ��  G� ��  J= ��  J= ��  G� ��  G�      D   , �C  @� �C  Cq �)  Cq �)  @� �C  @�      D   , �"  ;8 �"  <x �l  <x �l  ;8 �"  ;8      D   , �  K� �  L� �  L� �  K� �  K�      D   , �  G� �  J= �  J= �  G� �  G�      D   , ��  G� ��  I� �[  I� �[  G� ��  G�      D   , �  G� �  J= �  J= �  G� �  G�      D   , �  K� �  L� �  L� �  K� �  K�      D   , �  @� �  Cq �  Cq �  @� �  @�      D   , �  G� �  J= �  J= �  G� �  G�      D   , �  K� �  L� �  L� �  K� �  K�      D   , �  @� �  Cq �B  Cq �B  @� �  @�      D   , �  G� �  J= �  J= �  G� �  G�      D   , �  @� �  Cq �  Cq �  @� �  @�      D   , �  ;8 �  <x �B  <x �B  ;8 �  ;8      D   , �  K� �  L� �  L� �  K� �  K�      D   , �x  @� �x  Cq �  Cq �  @� �x  @�      D   , �  G� �  I� ��  I� ��  G� �  G�      D   , �/  @� �/  Cq �  Cq �  @� �/  @�      D   , �_  G� �_  I� ��  I� ��  G� �_  G�      D   , �  ;8 �  <x ��  <x ��  ;8 �  ;8      D   , ��  G� ��  I� �o  I� �o  G� ��  G�      D   , �_  G� �_  I� ��  I� ��  G� �_  G�      D   , �.  K� �.  L� �  L� �  K� �.  K�      D   , ��  @� ��  Cq ��  Cq ��  @� ��  @�      D   , �B  K� �B  L� ��  L� ��  K� �B  K�      D   , �/  G� �/  J= �  J= �  G� �/  G�      D   , �C  G� �C  J= �)  J= �)  G� �C  G�      D   , �/  @� �/  Cq �  Cq �  @� �/  @�      D   , ��  G� ��  J= ��  J= ��  G� ��  G�      D   , �  @� �  Cq ��  Cq ��  @� �  @�      D   , ��  G� ��  I� �3  I� �3  G� ��  G�      D   , �  >b �  ?p �n  ?p �n  >b �  >b      D   , �  K� �  L� �s  L� �s  K� �  K�      D   , ��  @� ��  Cq �  Cq �  @� ��  @�      D   , �  K� �  L� �x  L� �x  K� �  K�      D   , �  G� �  J= ��  J= ��  G� �  G�      D   , �N  >b �N  ?p َ  ?p َ  >b �N  >b      D   , �/  ;8 �/  <x �o  <x �o  ;8 �/  ;8      D   , �  %{ �  ,= ��  ,= ��  %{ �  %{      D   , ��   & ��  !� ��  !� ��   & ��   &      D   , ��   & ��  !� ��  !� ��   & ��   &      D   , �  # �  #� �x  #� �x  # �  #      D   , ��  '� ��  )� �3  )� �3  '� ��  '�      D   , �i  "� �i  $, ��  $, ��  "� �i  "�      D   , �  # �  #� �  #� �  # �  #      D   , ��   & ��  !� ��  !� ��   & ��   &      D   , �  "� �  $, �  $, �  "� �  "�      D   , ��  '� ��  )� �[  )� �[  '� ��  '�      D   , �   & �  !� �  !� �   & �   &      D   , �  0/ �  6� �  6� �  0/ �  0/      D   , �  %{ �  ,= �  ,= �  %{ �  %{      D   , �_  '� �_  )� ��  )� ��  '� �_  '�      D   , �  %{ �  ,= �  ,= �  %{ �  %{      D   , �_  '� �_  )� ��  )� ��  '� �_  '�      D   , �  %{ �  ,= �  ,= �  %{ �  %{      D   , �  %{ �  ,= �  ,= �  %{ �  %{      D   , ��   & ��  !� ��  !� ��   & ��   &      D   , �  # �  #� �  #� �  # �  #      D   , �  # �  #� �  #� �  # �  #      D   , �/  %{ �/  ,= �  ,= �  %{ �/  %{      D   , �C  %{ �C  ,= �)  ,= �)  %{ �C  %{      D   , ��  %{ ��  ,= ��  ,= ��  %{ ��  %{      D   , ��  0/ ��  6� ��  6� ��  0/ ��  0/      D   , �  # �  #� �*  #� �*  # �  #      D   , �/  0/ �/  6� �  6� �  0/ �/  0/      D   , ��  0/ ��  6� ��  6� ��  0/ ��  0/      D   , ��  '� ��  )� �o  )� �o  '� ��  '�      D   , �C  %{ �C  ,= �)  ,= �)  %{ �C  %{      D   , �.  "� �.  $, �  $, �  "� �.  "�      D   , �/  %{ �/  ,= �  ,= �  %{ �/  %{      D   , ��  %{ ��  ,= ��  ,= ��  %{ ��  %{      D   , �  0/ �  6� �  6� �  0/ �  0/      D   , �.  # �.  #� �  #� �  # �.  #      D   , �  0/ �  6� �B  6� �B  0/ �  0/      D   , ��  '� ��  )� �o  )� �o  '� ��  '�      D   , �  %{ �  ,= �  ,= �  %{ �  %{      D   , �  '� �  )� ��  )� ��  '� �  '�      D   , �B  # �B  #� ��  #� ��  # �B  #      D   , �  %{ �  ,= �  ,= �  %{ �  %{      D   , �   & �  !� 	�  !� 	�   & �   &      D   ,   K�   L� z  L� z  K�   K�      D   ,   K�   L� z  L� z  K�   K�      D   ,   #   #� z  #� z  #   #      D   ,   "�   $, z  $, z  "�   "�      D   , �  G� �  J= y  J= y  G� �  G�      D   , �  G� �  J= �  J= �  G� �  G�      D   , 
  K� 
  L� �  L� �  K� 
  K�      D   , �  ;8 �  <x F  <x F  ;8 �  ;8      D   , �  ;8 �  <x �  <x �  ;8 �  ;8      D   , z  ;8 z  <x �  <x �  ;8 z  ;8      D   , a  G� a  I� �  I� �  G� a  G�      D   , �  @� �  Cq �  Cq �  @� �  @�      D   , 1  G� 1  J=   J=   G� 1  G�      D   , 	  @� 	  Cq 
  Cq 
  @� 	  @�      D   , �  K� �  L�   L�   K� �  K�      D   , �  K� �  L� 	  L� 	  K� �  K�      D   , 0  K� 0  L� �  L� �  K� 0  K�      D   , �  @� �  Cq 
0  Cq 
0  @� �  @�      D   , �  K� �  L�   L�   K� �  K�      D   , 1  @� 1  Cq   Cq   @� 1  @�      D   , �  G� �  J= �  J= �  G� �  G�      D   , �  G� �  I� 
I  I� 
I  G� �  G�      D   , 	  G� 	  J= 
  J= 
  G� 	  G�      D   , �  @� �  Cq �  Cq �  @� �  @�      D   , �  G� �  I� 
I  I� 
I  G� �  G�      D   , u  G� u  I� �  I� �  G� u  G�      D   , 1  G� 1  J=   J=   G� 1  G�      D   , z  @� z  Cq �  Cq �  @� z  @�      D   , 	  G� 	  J= 
  J= 
  G� 	  G�      D   , �  G� �  J= �  J= �  G� �  G�      D   , ]  ;8 ]  <x �  <x �  ;8 ]  ;8      D   , 
&  >b 
&  ?p �  ?p �  >b 
&  >b      D   , �  G� �  J= y  J= y  G� �  G�      D   , �  @� �  Cq y  Cq y  @� �  @�      D   , ��  @� ��  Cq ��  Cq ��  @� ��  @�      D   , ��  G� ��  I� �  I� �  G� ��  G�      D   , �W  @� �W  Cq �=  Cq �=  @� �W  @�      D   , ��  G� ��  J= ��  J= ��  G� ��  G�      D   , �V  K� �V  L� ��  L� ��  K� �V  K�      D   , ��  ;8 ��  <x �
  <x �
  ;8 ��  ;8      D   , �W  G� �W  J= �=  J= �=  G� �W  G�      D   , ��  >b ��  ?p �H  ?p �H  >b ��  >b      D   , �^  ;8 �^  <x  �  <x  �  ;8 �^  ;8      D   , ��  G� ��  J= ��  J= ��  G� ��  G�      D   , �j  K� �j  L� ��  L� ��  K� �j  K�      D   ,   G�   J= e  J= e  G�   G�      D   , R  @� R  Cq �  Cq �  @� R  @�      D   , �W  G� �W  J= �=  J= �=  G� �W  G�      D   , �>  ;8 �>  <x �~  <x �~  ;8 �>  ;8      D   , �>  @� �>  Cq �~  Cq �~  @� �>  @�      D   , �  @� �  Cq   Cq   @� �  @�      D   , �k  G� �k  J= �Q  J= �Q  G� �k  G�      D   , 	  G� 	  J= �  J= �  G� 	  G�      D   , ��  @� ��  Cq ��  Cq ��  @� ��  @�      D   , �  G� �  I� 5  I� 5  G� �  G�      D   , �k  @� �k  Cq �Q  Cq �Q  @� �k  @�      D   ,   G�   J= e  J= e  G�   G�      D   , �k  @� �k  Cq �Q  Cq �Q  @� �k  @�      D   , 	  @� 	  Cq �  Cq �  @� 	  @�      D   , �%  G� �%  I� ��  I� ��  G� �%  G�      D   , ��  G� ��  J= ��  J= ��  G� ��  G�      D   , 9  G� 9  I� �  I� �  G� 9  G�      D   , ��  K� ��  L� �R  L� �R  K� ��  K�      D   , ~  K� ~  L� �  L� �  K� ~  K�      D   , �j  K� �j  L� ��  L� ��  K� �j  K�      D   , ��  G� ��  J= ��  J= ��  G� ��  G�      D   , �  ;8 �  <x   <x   ;8 �  ;8      D   , �k  G� �k  J= �Q  J= �Q  G� �k  G�      D   , 	  @� 	  Cq �  Cq �  @� 	  @�      D   , 	  G� 	  J= �  J= �  G� 	  G�      D   ,   @�   Cq e  Cq e  @�   @�      D   , 9  G� 9  I� �  I� �  G� 9  G�      D   , ��  K� ��  L� f  L� f  K� ��  K�      D   , ��  G� ��  I� �  I� �  G� ��  G�      D   , ��  @� ��  Cq ��  Cq ��  @� ��  @�      D   , �W  0/ �W  6� �=  6� �=  0/ �W  0/      D   , �V  # �V  #� ��  #� ��  # �V  #      D   , ��  %{ ��  ,= ��  ,= ��  %{ ��  %{      D   , �W  %{ �W  ,= �=  ,= �=  %{ �W  %{      D   , �/   & �/  !�    !�     & �/   &      D   , �W  %{ �W  ,= �=  ,= �=  %{ �W  %{      D   , ��  %{ ��  ,= ��  ,= ��  %{ ��  %{      D   , ��  '� ��  )� �  )� �  '� ��  '�      D   , �  0/ �  6�   6�   0/ �  0/      D   , ��  # ��  #� �R  #� �R  # ��  #      D   , �k  %{ �k  ,= �Q  ,= �Q  %{ �k  %{      D   , 	  %{ 	  ,= �  ,= �  %{ 	  %{      D   , ~  # ~  #� �  #� �  # ~  #      D   , �T   & �T  !� �  !� �   & �T   &      D   ,   %{   ,= e  ,= e  %{   %{      D   , �j  # �j  #� ��  #� ��  # �j  #      D   , �k  %{ �k  ,= �Q  ,= �Q  %{ �k  %{      D   , 	  %{ 	  ,= �  ,= �  %{ 	  %{      D   , 9  '� 9  )� �  )� �  '� 9  '�      D   , �/   & �/  !�    !�     & �/   &      D   , �%  '� �%  )� ��  )� ��  '� �%  '�      D   , �j  "� �j  $, ��  $, ��  "� �j  "�      D   , �k  0/ �k  6� �Q  6� �Q  0/ �k  0/      D   , 	  0/ 	  6� �  6� �  0/ 	  0/      D   , �>  0/ �>  6� �~  6� �~  0/ �>  0/      D   , ��  '� ��  )� �  )� �  '� ��  '�      D   , 9  '� 9  )� �  )� �  '� 9  '�      D   , ��  %{ ��  ,= ��  ,= ��  %{ ��  %{      D   , �  '� �  )� 5  )� 5  '� �  '�      D   , ��  %{ ��  ,= ��  ,= ��  %{ ��  %{      D   , ��  # ��  #� f  #� f  # ��  #      D   ,   %{   ,= e  ,= e  %{   %{      D   , ��  0/ ��  6� ��  6� ��  0/ ��  0/      D   , �  %{ �  ,= y  ,= y  %{ �  %{      D   , �  0/ �  6� y  6� y  0/ �  0/      D   , k   & k  !� S  !� S   & k   &      D   , �  %{ �  ,= y  ,= y  %{ �  %{      D   , k   & k  !� S  !� S   & k   &      D   , �  # �  #� 	  #� 	  # �  #      D   , �  '� �  )� 
I  )� 
I  '� �  '�      D   , �  %{ �  ,= �  ,= �  %{ �  %{      D   , 0  # 0  #� �  #� �  # 0  #      D   , 1  %{ 1  ,=   ,=   %{ 1  %{      D   , 	�   & 	�  !� .  !� .   & 	�   &      D   , 	  %{ 	  ,= 
  ,= 
  %{ 	  %{      D   , 1  0/ 1  6�   6�   0/ 1  0/      D   , z  0/ z  6� �  6� �  0/ z  0/      D   , �  # �  #�   #�   # �  #      D   , 
  # 
  #� �  #� �  # 
  #      D   , �  '� �  )� 
I  )� 
I  '� �  '�      D   , �  0/ �  6� �  6� �  0/ �  0/      D   , u  '� u  )� �  )� �  '� u  '�      D   , �  %{ �  ,= �  ,= �  %{ �  %{      D   , �  "� �  $,   $,   "� �  "�      D   , a  '� a  )� �  )� �  '� a  '�      D   , 	  %{ 	  ,= 
  ,= 
  %{ 	  %{      D   , 1  %{ 1  ,=   ,=   %{ 1  %{      D   , �  %{ �  ,= �  ,= �  %{ �  %{      E   , �  d� �  f:   f:   d� �  d�   	   E   !      �  N  g� N  [�   	   E   !      �  �  g� �  [�   	   E   !      �    W   [�   	   E   !      �  �  W& �  [�   	   E   !      �  �z  @� �z  I�   	   E   !      �  �  @� �  I�   	   E   !      �  �  @� �  I�   	   E   !      �  �T  @� �T  I�   	   E   !      �  �  @� �  I�   	   E   !      �  	�  @� 	�  I�   	   E   !     @  �  b� �  ;8   	   E   !     @  ��  b� ��  ;8   	   E   !       ��  _� ��  >b   	   E   !       �"  { �"  "�   	   E   !       ں  R0 ں  K�   	   E   !     @  ��  { ��  S�   	   E   !      �  �  \� �  S�   	   E   !      �  �T  \� �T  S�   	   E   !      �  �  \� �  S�   	   E   !      �  �  \� �  S�   	   E   !      �  	�  \� 	�  S�   	   E   !      �  �  o� �  [�   	   E   !      �  �  l� �  qH   	   E   !      �    l�   qH   	   E   !      �  �,  m� �,  Zs   	   E   !      �  ��  m� ��  Zs   	   E   !      �  �h  m� �h  Zs   	   E   !      �  �  0/ �  Cq   	   E   !      �  �  0/ �  Cq   	   E   !      �  �@  0/ �@  Cq   	   E   !      �  ��  0/ ��  Cq   	   E   !      �  |  0/ |  Cq   	   E   !      �    0/   Cq   	   E   !      �    m�   Zs   	   E   !      �  �  m� �  Zs      E   , �  N* �  O� �  O� �  N* �  N*      E   , ��  N* ��  O� �y  O� �y  N* ��  N*      E   , �U  N* �U  O� �=  O� �=  N* �U  N*      E   , ��  P� ��  R0 �>  R0 �>  P� ��  P�      E   , ��  y� ��  { �>  { �>  y� ��  y�      E   , ��  "� ��  $, �>  $, �>  "� ��  "�      E   , ��  K� ��  L� �>  L� �>  K� ��  K�      E   , k  |. k  }� S  }� S  |. k  |.      E   , �/  |. �/  }�    }�    |. �/  |.      E   , �/  |. �/  }�    }�    |. �/  |.      E   , k  p! k  qk S  qk S  p! k  p!      E   ,   W   X\ �  X\ �  W   W      E   , ��  S� ��  U� �  U� �  S� ��  S�      E   , ��  t ��  v �  v �  t ��  t      E   , ��  t ��  v �  v �  t ��  t      E   , ��  S� ��  U� �  U� �  S� ��  S�      E   , ��  Zs ��  \� ��  \� ��  Zs ��  Zs      E   , ��  al ��  b�    b�    al ��  al      E   , 9  S� 9  U� �  U� �  S� 9  S�      E   , f  al f  b� �  b� �  al f  al      E   , �  S� �  U� 
I  U� 
I  S� �  S�      E   , ��  f� ��  m�    m�    f� ��  f�      E   , 9  t 9  v �  v �  t 9  t      E   , f  f� f  m� �  m� �  f� f  f�      E   , �  t �  v 
I  v 
I  t �  t      E   , ��  Zs ��  \�    \�    Zs ��  Zs      E   , f  Zs f  \� �  \� �  Zs f  Zs      E   , 9  t 9  v �  v �  t 9  t      E   , ��  S� ��  U�  !  U�  !  S� ��  S�      E   , M  S� M  U� �  U� �  S� M  S�      E   , �j  P� �j  R0 ��  R0 ��  P� �j  P�      E   ,   P�   R0 z  R0 z  P�   P�      E   , 9  S� 9  U� �  U� �  S� 9  S�      E   , ��  t ��  v  !  v  !  t ��  t      E   , M  t M  v �  v �  t M  t      E   , *  [� *  \� j  \� j  [� *  [�      E   , 2  [� 2  \� r  \� r  [� 2  [�      E   , �  [� �  \� �  \� �  [� �  [�      E   , �  Z� �  [� ,  [� ,  Z� �  Z�      E   , p  Z� p  [� �  [� �  Z� p  Z�      E   , %  n� %  o� e  o� e  n� %  n�      E   , *  g *  h j  h j  g *  g      E   , �  l� �  m� ,  m� ,  l� �  l�      E   , p  l� p  m� �  m� �  l� p  l�      E   , �  e �  f �  f �  e �  e      E   , 2  e 2  f r  f r  e 2  e      E   , �  f� �  g� �  g� �  f� �  f�      E   , 2  f� 2  g� r  g� r  f� 2  f�      E   , -  d� -  f w  f w  d� -  d�      E   , �  d� �  f �  f �  d� �  d�      E   , -  f� -  g� w  g� w  f� -  f�      E   , �  f� �  g� �  g� �  f� �  f�      E   , R  Zs R  \� �  \� �  Zs R  Zs      E   , �  Zs �  \� 
0  \� 
0  Zs �  Zs      E   , �j  y� �j  { ��  { ��  y� �j  y�      E   ,   y�   { z  { z  y�   y�      E   , �  S� �  U� ��  U� ��  S� �  S�      E   , ]  al ]  b� �  b� �  al ]  al      E   , �*  al �*  b� �j  b� �j  al �*  al      E   , �  t �  v ��  v ��  t �  t      E   ,   W0   X> y  X> y  W0   W0      E   , �*  f� �*  m� �j  m� �j  f� �*  f�      E   , �*  Zs �*  \� �j  \� �j  Zs �*  Zs      E   , #  p? #  qM ~  qM ~  p? #  p?      E   , k  |. k  }� S  }� S  |. k  |.      E   , ��  |. ��  }� ��  }� ��  |. ��  |.      E   , �s  S� �s  U� ��  U� ��  S� �s  S�      E   , ��  |. ��  }� ��  }� ��  |. ��  |.      E   , �.  P� �.  R0 �  R0 �  P� �.  P�      E   , ��  |. ��  }� ��  }� ��  |. ��  |.      E   , ��  S� ��  U� �G  U� �G  S� ��  S�      E   , �_  S� �_  U� ��  U� ��  S� �_  S�      E   , ��  S� ��  U� �o  U� �o  S� ��  S�      E   , �  al �  b� ��  b� ��  al �  al      E   , ��  |. ��  }� ��  }� ��  |. ��  |.      E   , �  P� �  R0 �  R0 �  P� �  P�      E   , ��  S� ��  U� �3  U� �3  S� ��  S�      E   , �s  t �s  v ��  v ��  t �s  t      E   , �N  ^t �N  _� َ  _� َ  ^t �N  ^t      E   , �.  y� �.  { �  { �  y� �.  y�      E   , �5  S\ �5  T� ٧  T� ٧  S\ �5  S\      E   , ��  t ��  v �G  v �G  t ��  t      E   , �  P� �  R0 �  R0 �  P� �  P�      E   , �.  P� �.  R0 �  R0 �  P� �.  P�      E   , �  y� �  { �  { �  y� �  y�      E   , ��  S� ��  U� �o  U� �o  S� ��  S�      E   , ��  al ��  b� �.  b� �.  al ��  al      E   , �  f� �  m� ��  m� ��  f� �  f�      E   , �/  al �/  b� �o  b� �o  al �/  al      E   , �P  y� �P  { ��  { ��  y� �P  y�      E   , �_  S� �_  U� ��  U� ��  S� �_  S�      E   , ��  t ��  v �o  v �o  t ��  t      E   , �P  q� �P  xi �  xi �  q� �P  q�      E   , ��  f� ��  m� �.  m� �.  f� ��  f�      E   , �  Zs �  \� ��  \� ��  Zs �  Zs      E   , �i  y� �i  { ��  { ��  y� �i  y�      E   , �_  t �_  v ��  v ��  t �_  t      E   , �_  t �_  v ��  v ��  t �_  t      E   , ��  t ��  v �o  v �o  t ��  t      E   , �P  S� �P  V1 �  V1 �  S� �P  S�      E   , �x  Zs �x  \� �  \� �  Zs �x  Zs      E   , ��  Zs ��  \� �.  \� �.  Zs ��  Zs      E   , �  Zs �  \� �V  \� �V  Zs �  Zs      E   , ��  t ��  v �3  v �3  t ��  t      E   , �(  P� �(  R0 �  R0 �  P� �(  P�      E   , �  P� �  R0 �s  R0 �s  P� �  P�      E   , �i  "� �i  $, ��  $, ��  "� �i  "�      E   , �N  >b �N  ?p َ  ?p َ  >b �N  >b      E   , �  K� �  L� �s  L� �s  K� �  K�      E   , �/  ;8 �/  <x �o  <x �o  ;8 �/  ;8      E   , ��   & ��  !� ��  !� ��   & ��   &      E   , ��   & ��  !� ��  !� ��   & ��   &      E   , �_  '� �_  )� ��  )� ��  '� �_  '�      E   , ��  '� ��  )� �o  )� �o  '� ��  '�      E   , ��  0/ ��  6� ��  6� ��  0/ ��  0/      E   , �  "� �  $, �  $, �  "� �  "�      E   , �K  '� �K  )� �  )� �  '� �K  '�      E   , ��  '� ��  )� �[  )� �[  '� ��  '�      E   , �  '� �  )� ��  )� ��  '� �  '�      E   , �.  "� �.  $, �  $, �  "� �.  "�      E   , ��   & ��  !� ��  !� ��   & ��   &      E   , ��  ;8 ��  <x ��  <x ��  ;8 ��  ;8      E   , �d  ;8 �d  <x �  <x �  ;8 �d  ;8      E   , �_  '� �_  )� ��  )� ��  '� �_  '�      E   , ��  '� ��  )� �o  )� �o  '� ��  '�      E   , �  ;8 �  <x �B  <x �B  ;8 �  ;8      E   , �d  0/ �d  6� �  6� �  0/ �d  0/      E   , �  K� �  L� �  L� �  K� �  K�      E   , ��  G� ��  I� �3  I� �3  G� ��  G�      E   , �_  G� �_  I� ��  I� ��  G� �_  G�      E   , ��  G� ��  I� �o  I� �o  G� ��  G�      E   , �K  G� �K  I� �  I� �  G� �K  G�      E   , ��  G� ��  I� �[  I� �[  G� ��  G�      E   , �  G� �  I� ��  I� ��  G� �  G�      E   , �.  K� �.  L� �  L� �  K� �.  K�      E   , ��   & ��  !� ��  !� ��   & ��   &      E   , �  0/ �  6� �B  6� �B  0/ �  0/      E   , �d  @� �d  Cq �  Cq �  @� �d  @�      E   , �  @� �  Cq �B  Cq �B  @� �  @�      E   , �_  G� �_  I� ��  I� ��  G� �_  G�      E   , ��  G� ��  I� �o  I� �o  G� ��  G�      E   , ��  @� ��  Cq ��  Cq ��  @� ��  @�      E   , �  @� �  Cq �V  Cq �V  @� �  @�      E   , �x  @� �x  Cq �  Cq �  @� �x  @�      E   , ��  @� ��  Cq �  Cq �  @� ��  @�      E   , ��  '� ��  )� �3  )� �3  '� ��  '�      E   , ��  G� ��  I� �  I� �  G� ��  G�      E   , ]  ;8 ]  <x �  <x �  ;8 ]  ;8      E   , ��  '� ��  )� �  )� �  '� ��  '�      E   , k   & k  !� S  !� S   & k   &      E   , ��  '� ��  )� �  )� �  '� ��  '�      E   , k   & k  !� S  !� S   & k   &      E   , ��  G� ��  I� �  I� �  G� ��  G�      E   , �/   & �/  !�    !�     & �/   &      E   , ��  @� ��  Cq ��  Cq ��  @� ��  @�      E   , �/   & �/  !�    !�     & �/   &      E   , �>  ;8 �>  <x �~  <x �~  ;8 �>  ;8      E   , �%  '� �%  )� ��  )� ��  '� �%  '�      E   , �  '� �  )� 5  )� 5  '� �  '�      E   , a  '� a  )� �  )� �  '� a  '�      E   , �>  @� �>  Cq �~  Cq �~  @� �>  @�      E   , �j  "� �j  $, ��  $, ��  "� �j  "�      E   ,   "�   $, z  $, z  "�   "�      E   , �  "� �  $,   $,   "� �  "�      E   , �  @� �  Cq   Cq   @� �  @�      E   , �j  K� �j  L� ��  L� ��  K� �j  K�      E   , �%  G� �%  I� ��  I� ��  G� �%  G�      E   , �  G� �  I� 5  I� 5  G� �  G�      E   , a  G� a  I� �  I� �  G� a  G�      E   ,   K�   L� z  L� z  K�   K�      E   , 9  '� 9  )� �  )� �  '� 9  '�      E   , �  '� �  )� 
I  )� 
I  '� �  '�      E   , �  K� �  L�   L�   K� �  K�      E   , z  @� z  Cq �  Cq �  @� z  @�      E   , �  ;8 �  <x   <x   ;8 �  ;8      E   , �>  0/ �>  6� �~  6� �~  0/ �>  0/      E   , �  0/ �  6�   6�   0/ �  0/      E   , 9  G� 9  I� �  I� �  G� 9  G�      E   , �  G� �  I� 
I  I� 
I  G� �  G�      E   , u  G� u  I� �  I� �  G� u  G�      E   , z  0/ z  6� �  6� �  0/ z  0/      E   , 9  G� 9  I� �  I� �  G� 9  G�      E   , �  G� �  I� 
I  I� 
I  G� �  G�      E   , 9  '� 9  )� �  )� �  '� 9  '�      E   , �  '� �  )� 
I  )� 
I  '� �  '�      E   , u  '� u  )� �  )� �  '� u  '�      E   , z  ;8 z  <x �  <x �  ;8 z  ;8      E   , �  @� �  Cq 
0  Cq 
0  @� �  @�      E   , R  @� R  Cq �  Cq �  @� R  @�      D  , , �  e1 �  e� 1  e� 1  e1 �  e1      D  , , [  e1 [  e� �  e� �  e1 [  e1      D  , , 6  N� 6  O= �  O= �  N� 6  N�      D  , , ��  N� ��  O= ��  O= ��  N� ��  N�      D  , , �  N� �  O= �T  O= �T  N� �  N�      D  , , v  N� v  O=   O=   N� v  N�      D  , , �:  N� �:  O= ��  O= ��  N� �:  N�      D  , , ��  N� ��  O= �  O= �  N� ��  N�      D  , , �  N� �  O= L  O= L  N� �  N�      D  , , �z  N� �z  O= �  O= �  N� �z  N�      D  , , �>  N� �>  O= ��  O= ��  N� �>  N�      D  , , �  p{ �  q ^  q ^  p{ �  p{      D  , , �  |� �  }A j  }A j  |� �  |�      D  , , �  |� �  }A j  }A j  |� �  |�      D  , , ��  |� ��  }A �.  }A �.  |� ��  |�      D  , , ��  |� ��  }A �.  }A �.  |� ��  |�      D  , ,   Wl   X �  X �  Wl   Wl      D  , ,   p{   q �  q �  p{   p{      D  , , C  Wl C  X �  X �  Wl C  Wl      D  , ,   |�   }A �  }A �  |�   |�      D  , ,   |�   }A �  }A �  |�   |�      D  , , ��  |� ��  }A �n  }A �n  |� ��  |�      D  , , ��  |� ��  }A �n  }A �n  |� ��  |�      D  , , H  p{ H  q �  q �  p{ H  p{      D  , , �  a� �  bW H  bW H  a� �  a�      D  , , �  Wl �  X Y  X Y  Wl �  Wl      D  , , T  |� T  }A �  }A �  |� T  |�      D  , , T  |� T  }A �  }A �  |� T  |�      D  , , �  |� �  }A ��  }A ��  |� �  |�      D  , , �  |� �  }A ��  }A ��  |� �  |�      D  , , �  Z� �  [c =  [c =  Z� �  Z�      D  , , 	E  Z� 	E  [c 	�  [c 	�  Z� 	E  Z�      D  , , �	  Z� �	  [c ��  [c ��  Z� �	  Z�      D  , , �  \ �  \� =  \� =  \ �  \      D  , , 	E  \ 	E  \� 	�  \� 	�  \ 	E  \      D  , , �	  \ �	  \� ��  \� ��  \ �	  \      D  , ,   \!   \�   \�   \!   \!      D  , , �  \! �  \�   \�   \! �  \!      D  , ,   \!   \� �  \� �  \!   \!      D  , , A  Z� A  [O �  [O �  Z� A  Z�      D  , , �  Z� �  [O [  [O [  Z� �  Z�      D  , , z  n� z  oO   oO   n� z  n�      D  , ,   g9   g�   g�   g9   g9      D  , , A  l� A  mo �  mo �  l� A  l�      D  , , �  l� �  mo [  mo [  l� �  l�      D  , ,   e;   e� �  e� �  e;   e;      D  , , �  e; �  e�   e�   e; �  e;      D  , ,   g   g� �  g� �  g   g      D  , , �  g �  g�   g�   g �  g      D  , , �  e; �  e�   e�   e; �  e;      D  , ,   e;   e� �  e� �  e;   e;      D  , , �  g �  g�   g�   g �  g      D  , ,   g   g� �  g� �  g   g      D  , , �  a� �  bW ��  bW ��  a� �  a�      D  , , �  a� �  bW Q  bW Q  a� �  a�      D  , , �  g� �  h ��  h ��  g� �  g�      D  , , �  g� �  h Q  h Q  g� �  g�      D  , , �  h� �  i_ ��  i_ ��  h� �  h�      D  , , �  h� �  i_ Q  i_ Q  h� �  h�      D  , , �  j	 �  j� ��  j� ��  j	 �  j	      D  , , �  j	 �  j� Q  j� Q  j	 �  j	      D  , , �  kI �  k� ��  k� ��  kI �  kI      D  , , �  kI �  k� Q  k� Q  kI �  kI      D  , , �  l� �  m ��  m ��  l� �  l�      D  , , �  l� �  m Q  m Q  l� �  l�      D  , , �  Z� �  [c ��  [c ��  Z� �  Z�      D  , , �  Z� �  [c Q  [c Q  Z� �  Z�      D  , , �  \ �  \� ��  \� ��  \ �  \      D  , , �  \ �  \� Q  \� Q  \ �  \      D  , , ��  Q@ ��  Q� �n  Q� �n  Q@ ��  Q@      D  , , v  Q@ v  Q�   Q�   Q@ v  Q@      D  , , ��  z ��  z� �n  z� �n  z ��  z      D  , , v  z v  z�   z�   z v  z      D  , , �	  T� �	  U7 ��  U7 ��  T� �	  T�      D  , , �  T� �  U7 =  U7 =  T� �  T�      D  , , 	E  T� 	E  U7 	�  U7 	�  T� 	E  T�      D  , , �	  t� �	  uS ��  uS ��  t� �	  t�      D  , , �  t� �  uS =  uS =  t� �  t�      D  , , 	E  t� 	E  uS 	�  uS 	�  t� 	E  t�      D  , , �	  t� �	  uS ��  uS ��  t� �	  t�      D  , , �  t� �  uS =  uS =  t� �  t�      D  , , �  T� �  U7 ��  U7 ��  T� �  T�      D  , , �  T� �  U7 Q  U7 Q  T� �  T�      D  , , �	  T� �	  U7 ��  U7 ��  T� �	  T�      D  , , �  T� �  U7 =  U7 =  T� �  T�      D  , , �  t� �  uS ��  uS ��  t� �  t�      D  , , �  t� �  uS Q  uS Q  t� �  t�      D  , , �  l� �  m �  m �  l� �  l�      D  , , �  a� �  bW �  bW �  a� �  a�      D  , , �  Z� �  [c �  [c �  Z� �  Z�      D  , , �  \ �  \� �  \� �  \ �  \      D  , , �  g� �  h �  h �  g� �  g�      D  , , �:  Q@ �:  Q� ��  Q� ��  Q@ �:  Q@      D  , , �:  z �:  z� ��  z� ��  z �:  z      D  , , �  h� �  i_ �  i_ �  h� �  h�      D  , , �  j	 �  j� �  j� �  j	 �  j	      D  , , �  T� �  U7 �  U7 �  T� �  T�      D  , , �  kI �  k� �  k� �  kI �  kI      D  , , �  t� �  uS �  uS �  t� �  t�      D  , , ��  |� ��  }A �r  }A �r  |� ��  |�      D  , , ��  |� ��  }A �Z  }A �Z  |� ��  |�      D  , , ��  |� ��  }A �Z  }A �Z  |� ��  |�      D  , , أ  ^� أ  _F �9  _F �9  ^� أ  ^�      D  , , ��  z ��  z� �m  z� �m  z ��  z      D  , , �\  |� �\  }A ��  }A ��  |� �\  |�      D  , , ��  l� ��  m �w  m �w  l� ��  l�      D  , , �  |� �  }A �2  }A �2  |� �  |�      D  , , �  |� �  }A �2  }A �2  |� �  |�      D  , , �  s} �  t �;  t �;  s} �  s}      D  , , �C  l� �C  m ��  m ��  l� �C  l�      D  , , ��  Z� ��  [c �w  [c �w  Z� ��  Z�      D  , , ބ  |� ބ  }A �  }A �  |� ބ  |�      D  , , �  t� �  uS �;  uS �;  t� �  t�      D  , , �C  a� �C  bW ��  bW ��  a� �C  a�      D  , , �C  Z� �C  [c ��  [c ��  Z� �C  Z�      D  , , ��  \ ��  \� �w  \� �w  \ ��  \      D  , , ބ  |� ބ  }A �  }A �  |� ބ  |�      D  , , ��  g� ��  h �w  h �w  g� ��  g�      D  , , �\  |� �\  }A ��  }A ��  |� �\  |�      D  , , �C  \ �C  \� ��  \� ��  \ �C  \      D  , , �  Q@ �  Q� �2  Q� �2  Q@ �  Q@      D  , , �D  |� �D  }A ��  }A ��  |� �D  |�      D  , , �  u� �  v� �;  v� �;  u� �  u�      D  , , �  w= �  w� �;  w� �;  w= �  w=      D  , , ��  Q@ ��  Q� �  Q� �  Q@ ��  Q@      D  , , �  z �  z� �2  z� �2  z �  z      D  , , �D  |� �D  }A ��  }A ��  |� �D  |�      D  , , �C  g� �C  h ��  h ��  g� �C  g�      D  , , ��  h� ��  i_ �w  i_ �w  h� ��  h�      D  , , ��  z ��  z� �  z� �  z ��  z      D  , , �k  T� �k  U7 �  U7 �  T� �k  T�      D  , , ��  Q@ ��  Q� �,  Q� �,  Q@ ��  Q@      D  , , �k  Z� �k  [c �  [c �  Z� �k  Z�      D  , , �k  \ �k  \� �  \� �  \ �k  \      D  , , ��  T� ��  U7 �c  U7 �c  T� ��  T�      D  , , �k  t� �k  uS �  uS �  t� �k  t�      D  , , �C  h� �C  i_ ��  i_ ��  h� �C  h�      D  , , ��  j	 ��  j� �w  j� �w  j	 ��  j	      D  , , �o  Q@ �o  Q� �  Q� �  Q@ �o  Q@      D  , , ��  t� ��  uS �c  uS �c  t� ��  t�      D  , , ��  t� ��  uS �c  uS �c  t� ��  t�      D  , , �k  t� �k  uS �  uS �  t� �k  t�      D  , , �  r= �  r� �;  r� �;  r= �  r=      D  , , ��  Q@ ��  Q� �  Q� �  Q@ ��  Q@      D  , , �/  t� �/  uS ��  uS ��  t� �/  t�      D  , , ��  T� ��  U7 �w  U7 �w  T� ��  T�      D  , , أ  S� أ  TL �9  TL �9  S� أ  S�      D  , , �C  j	 �C  j� ��  j� ��  j	 �C  j	      D  , , ��  kI ��  k� �w  k� �w  kI ��  kI      D  , , �C  T� �C  U7 ��  U7 ��  T� �C  T�      D  , , ��  T� ��  U7 �c  U7 �c  T� ��  T�      D  , , �k  T� �k  U7 �  U7 �  T� �k  T�      D  , , ބ  a� ބ  bW �  bW �  a� ބ  a�      D  , , �  Q@ �  Q� �2  Q� �2  Q@ �  Q@      D  , , �/  T� �/  U7 ��  U7 ��  T� �/  T�      D  , , ��  t� ��  uS �w  uS �w  t� ��  t�      D  , , ��  |� ��  }A �r  }A �r  |� ��  |�      D  , , ��  a� ��  bW �w  bW �w  a� ��  a�      D  , , �C  kI �C  k� ��  k� ��  kI �C  kI      D  , , �C  t� �C  uS ��  uS ��  t� �C  t�      D  , , �  z �  z� �J  z� �J  z �  z      D  , , ��  z ��  z� �  z� �  z ��  z      D  , , �  T �  T� �;  T� �;  T �  T      D  , , ��  Z� ��  [c �c  [c �c  Z� ��  Z�      D  , , �  UA �  U� �;  U� �;  UA �  UA      D  , , ��  \ ��  \� �c  \� �c  \ ��  \      D  , , أ  >� أ  ?4 �9  ?4 �9  >� أ  >�      D  , , ��  #< ��  #� �m  #� �m  #< ��  #<      D  , , �o  L �o  L� �  L� �  L �o  L      D  , , �   � �  !9 �2  !9 �2   � �   �      D  , , �   � �  !9 �2  !9 �2   � �   �      D  , , ބ   � ބ  !9 �  !9 �   � ބ   �      D  , , ��   � ��  !9 �r  !9 �r   � ��   �      D  , , ��   � ��  !9 �r  !9 �r   � ��   �      D  , , ��   � ��  !9 �Z  !9 �Z   � ��   �      D  , , ��   � ��  !9 �Z  !9 �Z   � ��   �      D  , , ބ   � ބ  !9 �  !9 �   � ބ   �      D  , , ބ  ;� ބ  <# �  <# �  ;� ބ  ;�      D  , , �\   � �\  !9 ��  !9 ��   � �\   �      D  , , �\   � �\  !9 ��  !9 ��   � �\   �      D  , , �D   � �D  !9 ��  !9 ��   � �D   �      D  , , �D   � �D  !9 ��  !9 ��   � �D   �      D  , , �W  0� �W  1[ ��  1[ ��  0� �W  0�      D  , , ��  0� ��  1[ ��  1[ ��  0� ��  0�      D  , , ��  AA ��  A� �c  A� �c  AA ��  AA      D  , , �/  H� �/  IC ��  IC ��  H� �/  H�      D  , , ��  H� ��  IC �c  IC �c  H� ��  H�      D  , , �k  H� �k  IC �  IC �  H� �k  H�      D  , , �/  AA �/  A� ��  A� ��  AA �/  AA      D  , , ��  B� ��  C �c  C �c  B� ��  B�      D  , , �/  B� �/  C ��  C ��  B� �/  B�      D  , , �  5� �  6[ �O  6[ �O  5� �  5�      D  , , �  B� �  C �O  C �O  B� �  B�      D  , , �/  (� �/  )' ��  )' ��  (� �/  (�      D  , , ��  (� ��  )' �c  )' �c  (� ��  (�      D  , , �k  (� �k  )' �  )' �  (� �k  (�      D  , , �W  B� �W  C ��  C ��  B� �W  B�      D  , , ��  B� ��  C ��  C ��  B� ��  B�      D  , , �  3E �  3� �O  3� �O  3E �  3E      D  , , �W  3E �W  3� ��  3� ��  3E �W  3E      D  , , ��  3E ��  3� ��  3� ��  3E ��  3E      D  , , ��  (� ��  )' �c  )' �c  (� ��  (�      D  , , �k  (� �k  )' �  )' �  (� �k  (�      D  , , �W  5� �W  6[ ��  6[ ��  5� �W  5�      D  , , ��  5� ��  6[ ��  6[ ��  5� ��  5�      D  , , �  AA �  A� �O  A� �O  AA �  AA      D  , , �W  AA �W  A� ��  A� ��  AA �W  AA      D  , , ��  AA ��  A� ��  A� ��  AA ��  AA      D  , , �  H� �  IC �O  IC �O  H� �  H�      D  , , �W  H� �W  IC ��  IC ��  H� �W  H�      D  , , ��  H� ��  IC ��  IC ��  H� ��  H�      D  , , �k  B� �k  C �  C �  B� �k  B�      D  , , �  ;� �  <# �O  <# �O  ;� �  ;�      D  , , �W  ;� �W  <# ��  <# ��  ;� �W  ;�      D  , , �  2 �  2� �O  2� �O  2 �  2      D  , , �W  2 �W  2� ��  2� ��  2 �W  2      D  , , ��  H� ��  IC �c  IC �c  H� ��  H�      D  , , �k  H� �k  IC �  IC �  H� �k  H�      D  , , ��  L ��  L� �  L� �  L ��  L      D  , , �  L �  L� �2  L� �2  L �  L      D  , , ��  2 ��  2� ��  2� ��  2 ��  2      D  , , ��  ;� ��  <# ��  <# ��  ;� ��  ;�      D  , , �  (� �  )' �O  )' �O  (� �  (�      D  , , �W  (� �W  )' ��  )' ��  (� �W  (�      D  , , ��  (� ��  )' ��  )' ��  (� ��  (�      D  , , �k  AA �k  A� �  A� �  AA �k  AA      D  , , �  4� �  5 �O  5 �O  4� �  4�      D  , , �W  4� �W  5 ��  5 ��  4� �W  4�      D  , , ��  #< ��  #� �  #� �  #< ��  #<      D  , , �  #< �  #� �2  #� �2  #< �  #<      D  , , ��  4� ��  5 ��  5 ��  4� ��  4�      D  , , �  0� �  1[ �O  1[ �O  0� �  0�      D  , , �   � �  !9 ��  !9 ��   � �   �      D  , , �:  L �:  L� ��  L� ��  L �:  L      D  , ,    �   !9 �  !9 �   �    �      D  , , ��   � ��  !9 �n  !9 �n   � ��   �      D  , , ��   � ��  !9 �n  !9 �n   � ��   �      D  , , �  ;� �  <# H  <# H  ;� �  ;�      D  , , �   � �  !9 j  !9 j   � �   �      D  , , �   � �  !9 j  !9 j   � �   �      D  , , ��   � ��  !9 �.  !9 �.   � ��   �      D  , , ��   � ��  !9 �.  !9 �.   � ��   �      D  , ,    �   !9 �  !9 �   �    �      D  , , T   � T  !9 �  !9 �   � T   �      D  , , �:  #< �:  #� ��  #� ��  #< �:  #<      D  , , T   � T  !9 �  !9 �   � T   �      D  , , �   � �  !9 ��  !9 ��   � �   �      D  , , 	E  B� 	E  C 	�  C 	�  B� 	E  B�      D  , , �	  (� �	  )' ��  )' ��  (� �	  (�      D  , , �  (� �  )' =  )' =  (� �  (�      D  , , 	E  (� 	E  )' 	�  )' 	�  (� 	E  (�      D  , , �  B� �  C =  C =  B� �  B�      D  , , �	  B� �	  C ��  C ��  B� �	  B�      D  , , ��  3E ��  3� �)  3� �)  3E ��  3E      D  , , ��  0� ��  1[ �)  1[ �)  0� ��  0�      D  , , 1  0� 1  1[ �  1[ �  0� 1  0�      D  , , �  0� �  1[ e  1[ e  0� �  0�      D  , , ��  L ��  L� �n  L� �n  L ��  L      D  , , �	  (� �	  )' ��  )' ��  (� �	  (�      D  , , �  (� �  )' =  )' =  (� �  (�      D  , , 	E  (� 	E  )' 	�  )' 	�  (� 	E  (�      D  , , �  (� �  )' y  )' y  (� �  (�      D  , , v  L v  L�   L�   L v  L      D  , ,   L   L� �  L� �  L   L      D  , , 1  3E 1  3� �  3� �  3E 1  3E      D  , , �  3E �  3� e  3� e  3E �  3E      D  , , �	  AA �	  A� ��  A� ��  AA �	  AA      D  , , 	E  AA 	E  A� 	�  A� 	�  AA 	E  AA      D  , , �  AA �  A� =  A� =  AA �  AA      D  , , ��  ;� ��  <# �)  <# �)  ;� ��  ;�      D  , , ��  H� ��  IC �)  IC �)  H� ��  H�      D  , , 1  H� 1  IC �  IC �  H� 1  H�      D  , , �  H� �  IC e  IC e  H� �  H�      D  , , ��  4� ��  5 �)  5 �)  4� ��  4�      D  , , 1  4� 1  5 �  5 �  4� 1  4�      D  , , ��  #< ��  #� �n  #� �n  #< ��  #<      D  , , v  #< v  #�   #�   #< v  #<      D  , ,   #<   #� �  #� �  #<   #<      D  , , ��  B� ��  C �)  C �)  B� ��  B�      D  , , 1  B� 1  C �  C �  B� 1  B�      D  , , �	  H� �	  IC ��  IC ��  H� �	  H�      D  , , �  H� �  IC =  IC =  H� �  H�      D  , , 	E  H� 	E  IC 	�  IC 	�  H� 	E  H�      D  , , �  H� �  IC y  IC y  H� �  H�      D  , , �  B� �  C e  C e  B� �  B�      D  , , �  4� �  5 e  5 e  4� �  4�      D  , , 1  ;� 1  <# �  <# �  ;� 1  ;�      D  , , ��  2 ��  2� �)  2� �)  2 ��  2      D  , , 1  2 1  2� �  2� �  2 1  2      D  , , �  2 �  2� e  2� e  2 �  2      D  , , �	  H� �	  IC ��  IC ��  H� �	  H�      D  , , �  H� �  IC =  IC =  H� �  H�      D  , , ��  (� ��  )' �)  )' �)  (� ��  (�      D  , , 1  (� 1  )' �  )' �  (� 1  (�      D  , , �  (� �  )' e  )' e  (� �  (�      D  , , 	E  H� 	E  IC 	�  IC 	�  H� 	E  H�      D  , , ��  5� ��  6[ �)  6[ �)  5� ��  5�      D  , , 1  5� 1  6[ �  6[ �  5� 1  5�      D  , , �  5� �  6[ e  6[ e  5� �  5�      D  , , ��  AA ��  A� �)  A� �)  AA ��  AA      D  , , 1  AA 1  A� �  A� �  AA 1  AA      D  , , �  AA �  A� e  A� e  AA �  AA      D  , , �  ;� �  <# e  <# e  ;� �  ;�      E  , , �  e �  e� r  e� r  e �  e      E  , ,   e   e� �  e� �  e   e      E  , , �  N� �  OV ]  OV ]  N� �  N�      E  , , �Y  N� �Y  OV �!  OV �!  N� �Y  N�      E  , , �  N� �  OV ��  OV ��  N� �  N�      E  , , %  N� %  OV �  OV �  N� %  N�      E  , , ��  N� ��  OV ��  OV ��  N� ��  N�      E  , , �  N� �  OV �u  OV �u  N� �  N�      E  , , ��  H� ��  I\ ��  I\ ��  H� ��  H�      E  , , ��  (x ��  )@ ��  )@ ��  (x ��  (x      E  , , 3  |� 3  }Z �  }Z �  |� 3  |�      E  , , ��  |� ��  }Z ��  }Z ��  |� ��  |�      E  , , �  |� �  }Z �  }Z �  |� �  |�      E  , , �  |� �  }Z �  }Z �  |� �  |�      E  , , ��  |� ��  }Z �O  }Z �O  |� ��  |�      E  , , ��  |� ��  }Z �O  }Z �O  |� ��  |�      E  , , �  WS �  X �  X �  WS �  WS      E  , , �  WS �  X T  X T  WS �  WS      E  , , 3  pb 3  q* �  q* �  pb 3  pb      E  , , �  pb �  q* �  q* �  pb �  pb      E  , , �!  Q' �!  Q� ��  Q� ��  Q' �!  Q'      E  , , ��  Q' ��  Q� ��  Q� ��  Q' ��  Q'      E  , , ]  Q' ]  Q� %  Q� %  Q' ]  Q'      E  , , �!  y� �!  z� ��  z� ��  y� �!  y�      E  , , ��  y� ��  z� ��  z� ��  y� ��  y�      E  , , ]  y� ]  z� %  z� %  y� ]  y�      E  , , ��  T� ��  UP ��  UP ��  T� ��  T�      E  , , �  T� �  UP V  UP V  T� �  T�      E  , , 	,  T� 	,  UP 	�  UP 	�  T� 	,  T�      E  , , ��  t� ��  ul ��  ul ��  t� ��  t�      E  , , �  t� �  ul V  ul V  t� �  t�      E  , , 	,  t� 	,  ul 	�  ul 	�  t� 	,  t�      E  , , ��  t� ��  ul ��  ul ��  t� ��  t�      E  , , �  t� �  ul V  ul V  t� �  t�      E  , , �f  T� �f  UP �.  UP �.  T� �f  T�      E  , , �  T� �  UP ��  UP ��  T� �  T�      E  , , ��  |� ��  }Z ��  }Z ��  |� ��  |�      E  , , �  T� �  UP j  UP j  T� �  T�      E  , , ��  T� ��  UP ��  UP ��  T� ��  T�      E  , , �  T� �  UP V  UP V  T� �  T�      E  , , �f  t� �f  ul �.  ul �.  t� �f  t�      E  , , �  t� �  ul ��  ul ��  t� �  t�      E  , , 3  |� 3  }Z �  }Z �  |� 3  |�      E  , , �  t� �  ul j  ul j  t� �  t�      E  , , ��  y� ��  z� �  z� �  y� ��  y�      E  , , �R  T� �R  UP �  UP �  T� �R  T�      E  , , �V  Q' �V  Q� �  Q� �  Q' �V  Q'      E  , , ؊  S� ؊  Te �R  Te �R  S� ؊  S�      E  , , ݣ  |� ݣ  }Z �k  }Z �k  |� ݣ  |�      E  , , �  T� �  UP �|  UP �|  T� �  T�      E  , , �R  t� �R  ul �  ul �  t� �R  t�      E  , , �  |� �  }Z �  }Z �  |� �  |�      E  , , �  |� �  }Z �  }Z �  |� �  |�      E  , , ݣ  |� ݣ  }Z �k  }Z �k  |� ݣ  |�      E  , , �  t� �  ul �|  ul �|  t� �  t�      E  , , �  t� �  ul �|  ul �|  t� �  t�      E  , , �R  t� �R  ul �  ul �  t� �R  t�      E  , , ��  Q' ��  Q� �  Q� �  Q' ��  Q'      E  , , �  Q' �  Q� �K  Q� �K  Q' �  Q'      E  , , �  t� �  ul ��  ul ��  t� �  t�      E  , , ��  T� ��  UP �  UP �  T� ��  T�      E  , , �;  y� �;  z� �  z� �  y� �;  y�      E  , , �  Q' �  Q� �K  Q� �K  Q' �  Q'      E  , , �K  |� �K  }Z �  }Z �  |� �K  |�      E  , , �K  |� �K  }Z �  }Z �  |� �K  |�      E  , , �*  T� �*  UP ��  UP ��  T� �*  T�      E  , , �  T� �  UP �|  UP �|  T� �  T�      E  , , �R  T� �R  UP �  UP �  T� �R  T�      E  , , �3  |� �3  }Z ��  }Z ��  |� �3  |�      E  , , ��  Q' ��  Q� �  Q� �  Q' ��  Q'      E  , , �  T� �  UP ��  UP ��  T� �  T�      E  , , ��  t� ��  ul �  ul �  t� ��  t�      E  , , �  y� �  z� �K  z� �K  y� �  y�      E  , , �3  |� �3  }Z ��  }Z ��  |� �3  |�      E  , , ־  y� ־  z� ׆  z� ׆  y� ־  y�      E  , , �}  Q' �}  Q� �E  Q� �E  Q' �}  Q'      E  , , �*  t� �*  ul ��  ul ��  t� �*  t�      E  , , �   � �  !R �  !R �   � �   �      E  , , �  (x �  )@ �|  )@ �|  (x �  (x      E  , , �R  (x �R  )@ �  )@ �  (x �R  (x      E  , , �   � �  !R �  !R �   � �   �      E  , , ݣ   � ݣ  !R �k  !R �k   � ݣ   �      E  , , ־  ## ־  #� ׆  #� ׆  ## ־  ##      E  , , �V  K� �V  L� �  L� �  K� �V  K�      E  , , �  H� �  I\ ��  I\ ��  H� �  H�      E  , , �  H� �  I\ �h  I\ �h  H� �  H�      E  , , �>  H� �>  I\ �  I\ �  H� �>  H�      E  , , �  H� �  I\ �|  I\ �|  H� �  H�      E  , , �R  H� �R  I\ �  I\ �  H� �R  H�      E  , , ��  K� ��  L� �  L� �  K� ��  K�      E  , , �  K� �  L� �K  L� �K  K� �  K�      E  , , �K   � �K  !R �  !R �   � �K   �      E  , , �K   � �K  !R �  !R �   � �K   �      E  , , �  H� �  I\ �|  I\ �|  H� �  H�      E  , , �R  H� �R  I\ �  I\ �  H� �R  H�      E  , , �3   � �3  !R ��  !R ��   � �3   �      E  , , �  (x �  )@ ��  )@ ��  (x �  (x      E  , , �  (x �  )@ �|  )@ �|  (x �  (x      E  , , �R  (x �R  )@ �  )@ �  (x �R  (x      E  , , �3   � �3  !R ��  !R ��   � �3   �      E  , , �  (x �  )@ �h  )@ �h  (x �  (x      E  , , �>  (x �>  )@ �  )@ �  (x �>  (x      E  , , ݣ   � ݣ  !R �k  !R �k   � ݣ   �      E  , , ��  ## ��  #� �  #� �  ## ��  ##      E  , , �  ## �  #� �K  #� �K  ## �  ##      E  , , �  (x �  )@ �  )@ �  (x �  (x      E  , , �   � �  !R �  !R �   � �   �      E  , , ��  H� ��  I\ ��  I\ ��  H� ��  H�      E  , , �  H� �  I\ V  I\ V  H� �  H�      E  , , 	,  H� 	,  I\ 	�  I\ 	�  H� 	,  H�      E  , , �   � �  !R �  !R �   � �   �      E  , , ��   � ��  !R �O  !R �O   � ��   �      E  , , ��   � ��  !R �O  !R �O   � ��   �      E  , , ��   � ��  !R ��  !R ��   � ��   �      E  , , �z  H� �z  I\ �B  I\ �B  H� �z  H�      E  , ,   H�   I\ �  I\ �  H�   H�      E  , , �  H� �  I\ ~  I\ ~  H� �  H�      E  , , �!  ## �!  #� ��  #� ��  ## �!  ##      E  , , ��  ## ��  #� ��  #� ��  ## ��  ##      E  , , ]  ## ]  #� %  #� %  ## ]  ##      E  , , �  ## �  #� �  #� �  ## �  ##      E  , , ��  (x ��  )@ ��  )@ ��  (x ��  (x      E  , , �  (x �  )@ V  )@ V  (x �  (x      E  , , 	,  (x 	,  )@ 	�  )@ 	�  (x 	,  (x      E  , , ��  H� ��  I\ ��  I\ ��  H� ��  H�      E  , , �  H� �  I\ V  I\ V  H� �  H�      E  , , 	,  H� 	,  I\ 	�  I\ 	�  H� 	,  H�      E  , , �  H� �  I\ �  I\ �  H� �  H�      E  , , 3   � 3  !R �  !R �   � 3   �      E  , , �!  K� �!  L� ��  L� ��  K� �!  K�      E  , , ��  K� ��  L� ��  L� ��  K� ��  K�      E  , , ]  K� ]  L� %  L� %  K� ]  K�      E  , , �  K� �  L� �  L� �  K� �  K�      E  , , 3   � 3  !R �  !R �   � 3   �      E  , , ��   � ��  !R ��  !R ��   � ��   �      E  , , ��  (x ��  )@ ��  )@ ��  (x ��  (x      E  , , �z  (x �z  )@ �B  )@ �B  (x �z  (x      E  , ,   (x   )@ �  )@ �  (x   (x      E  , , �  (x �  )@ ~  )@ ~  (x �  (x      E  , , �  (x �  )@ V  )@ V  (x �  (x      E  , , 	,  (x 	,  )@ 	�  )@ 	�  (x 	,  (x      �   ,             q� t� q� t�                  G      �"  |. vss       G      �  | vss       G        @L������ BZ        2l o� clk       G        @L������ BZ        =4 o� ena       G        @L������ BZ        '� o� 
rst_n       G        @�������  R�  � 
ua[0]       G        @�������  L  � 
ua[1]       G        @�������  ��  � 
ua[2]       G        @�������  p\  � 
ua[3]       G        @�������  $�  � 
ua[4]       G        @�������   �l  � 
ua[5]       G        @�������   ��  � 
ua[6]       G        @�������   B|  � 
ua[7]       G        @L������ BZ        � o� ui_in[0]      G        @L������ BZ         o� ui_in[1]      G        @L������ BZ        L o� ui_in[2]      G        @L������ BZ        �� o� ui_in[3]      G        @L������ BZ        � o� ui_in[4]      G        @L������ BZ        �� o� ui_in[5]      G        @L������ BZ        �, o� ui_in[6]      G        @L������ BZ        �d o� ui_in[7]      G        @L������ BZ        Ɯ o� uio_in[0]       G        @L������ BZ        �� o� uio_in[1]       G        @L������ BZ        � o� uio_in[2]       G        @L������ BZ        �D o� uio_in[3]       G        @L������ BZ        �| o� uio_in[4]       G        @L������ BZ        �� o� uio_in[5]       G        @L������ BZ        �� o� uio_in[6]       G        @L������ BZ        {$ o� uio_in[7]       G        @L������ BZ         �� o� uio_oe[0]       G        @L������ BZ         � o� uio_oe[1]       G        @L������ BZ         �L o� uio_oe[2]       G        @L������ BZ         �� o� uio_oe[3]       G        @L������ BZ         �� o� uio_oe[4]       G        @L������ BZ         �� o� uio_oe[5]       G        @L������ BZ         �, o� uio_oe[6]       G        @L������ BZ         xd o� uio_oe[7]       G        @L������ BZ         o� uio_out[0]      G        @L������ BZ        T o� uio_out[1]      G        @L������ BZ        � o� uio_out[2]      G        @L������ BZ         �� o� uio_out[3]      G        @L������ BZ         �� o� uio_out[4]      G        @L������ BZ         �4 o� uio_out[5]      G        @L������ BZ         �l o� uio_out[6]      G        @L������ BZ         Τ o� uio_out[7]      G        @L������ BZ        p\ o� uo_out[0]       G        @L������ BZ        e� o� uo_out[1]       G        @L������ BZ        Z� o� uo_out[2]       G        @L������ BZ        P o� uo_out[3]       G        @L������ BZ        E< o� uo_out[4]       G        @L������ BZ        :t o� uo_out[5]       G        @L������ BZ        /� o� uo_out[6]       G        @L������ BZ        $� o� uo_out[7]       G    	    @@         � �� 
VDPWR       G    	    @@         � �� VGND      G   , 1� m� 1� q� 3 q� 3 m� 1� m�      G   , <� m� <� q� =� q� =� m� <� m�      G   , ' m� ' q� (: q� (: m� ' m�      G   , Q     Q  � T�  � T�     Q          G   , �     �  � 	  � 	     �          G   , �     �  � ��  � ��     �          G   , n�     n�  � r  � r     n�          G   , #"     #"  � &�  � &�     #"          G   ,  ת      ת  �  �.  �  �.      ת          G   ,  �2      �2  �  ��  �  ��      �2          G   ,  @�      @�  �  D>  �  D>      @�          G   , F m� F q� r q� r m� F m�      G   , ~ m� ~ q� � q� � m� ~ m�      G   , � m� � q� � q� � m� � m�      G   , �� m� �� q� � q� � m� �� m�      G   , �& m� �& q� �R q� �R m� �& m�      G   , �^ m� �^ q� � q� � m� �^ m�      G   , ۖ m� ۖ q� �� q� �� m� ۖ m�      G   , �� m� �� q� �� q� �� m� �� m�      G   , � m� � q� �2 q� �2 m� � m�      G   , �> m� �> q� �j q� �j m� �> m�      G   , �v m� �v q� �� q� �� m� �v m�      G   , �� m� �� q� �� q� �� m� �� m�      G   , �� m� �� q� � q� � m� �� m�      G   , � m� � q� �J q� �J m� � m�      G   , �V m� �V q� �� q� �� m� �V m�      G   , z� m� z� q� {� q� {� m� z� m�      G   ,  �F m�  �F q�  �r q�  �r m�  �F m�      G   ,  �~ m�  �~ q�  �� q�  �� m�  �~ m�      G   ,  �� m�  �� q�  �� q�  �� m�  �� m�      G   ,  �� m�  �� q�  � q�  � m�  �� m�      G   ,  �& m�  �& q�  �R q�  �R m�  �& m�      G   ,  �^ m�  �^ q�  �� q�  �� m�  �^ m�      G   ,  �� m�  �� q�  �� q�  �� m�  �� m�      G   ,  w� m�  w� q�  x� q�  x� m�  w� m�      G   , � m� � q� � q� � m� � m�      G   , � m� � q� � q� � m� � m�      G   , � m� � q� " q� " m� � m�      G   ,  �. m�  �. q�  �Z q�  �Z m�  �. m�      G   ,  �f m�  �f q�  � q�  � m�  �f m�      G   ,  � m�  � q�  �� q�  �� m�  � m�      G   ,  �� m�  �� q�  � q�  � m�  �� m�      G   ,  � m�  � q�  �: q�  �: m�  � m�      G   , o� m� o� q� p� q� p� m� o� m�      G   , d� m� d� q� f* q� f* m� d� m�      G   , Z6 m� Z6 q� [b q� [b m� Z6 m�      G   , On m� On q� P� q� P� m� On m�      G   , D� m� D� q� E� q� E� m� D� m�      G   , 9� m� 9� q� ;
 q� ;
 m� 9� m�      G   , / m� / q� 0B q� 0B m� / m�      G   , $N m� $N q� %z q� %z m� $N m�      G   ,  �  �  � ^X  � ^X  �  �  �  �      G   ,  �  �  � ^X  p ^X  p  �  �  �      G      �"  |� vss       G      �  |� vss       A  , , �F  |. �F  }� ��  }� ��  |. �F  |.      A  , , ��  |. ��  }� �z  }� �z  |. ��  |.      A  , , �  W& �  XH �  XH �  W& �  W&      A  , , �  p5 �  qW �  qW �  p5 �  p5      A  , , ��  N* ��  O� �z  O� �z  N* ��  N*      A  , , �F  N* �F  O� ��  O� ��  N* �F  N*      A  , , �  |. �  }� �  }� �  |. �  |.      A  , , �  |. �  }� �T  }� �T  |. �  |.      A  , , �T  |. �T  }� �  }� �  |. �T  |.      A  , , �z   & �z  !� �  !� �   & �z   &      A  , , �   & �  !� �  !� �   & �   &      A  , , �   & �  !� �T  !� �T   & �   &      A  , , �T   & �T  !� �  !� �   & �T   &      A  , , �   & �  !� 	�  !� 	�   & �   &      A  , , 	�   & 	�  !� .  !� .   & 	�   &      A  , , �  |. �  }� 	�  }� 	�  |. �  |.      A  , , �z  |. �z  }� �  }� �  |. �z  |.      A  , , �  N* �  O� �  O� �  N* �  N*      A  , , �  N* �  O� �T  O� �T  N* �  N*      A  , , �T  N* �T  O� �  O� �  N* �T  N*      A  , , �z  N* �z  O� �  O� �  N* �z  N*      A  , , �  N* �  O� �  O� �  N* �  N*      A  , , �  N* �  O� �T  O� �T  N* �  N*      A  , , �T  N* �T  O� �  O� �  N* �T  N*      A  , , �  N* �  O� 	�  O� 	�  N* �  N*      A  , , 	�  N* 	�  O� .  O� .  N* 	�  N*      A  , , �  N* �  O� 	�  O� 	�  N* �  N*      A  , , �z  N* �z  O� �  O� �  N* �z  N*      ]  , , ��  {� ��  ~; �]  ~; �]  {� ��  {�      ]  , , �c  {� �c  ~; ��  ~; ��  {� �c  {�      ]  , , o  o� o  q�   q�   o� o  o�      ]  , , �  YG �  ^) �?  ^) �?  YG �  YG      ]  , , �-  YG �-  ^) ��  ^) ��  YG �-  YG      ]  , , ��  YG ��  ^)  {  ^)  {  YG ��  YG      ]  , , ��  ?� ��  D� �  D� �  ?� ��  ?�      ]  , , �  ?� �  D� �?  D� �?  ?� �  ?�      ]  , , �-  ?� �-  D� ��  D� ��  ?� �-  ?�      ]  , , ��  ?� ��  D�  {  D�  {  ?� ��  ?�      ]  , , i  ?� i  D�   D�   ?� i  ?�      ]  , ,   ?�   D� �  D� �  ?�   ?�      ]  , , i  YG i  ^)   ^)   YG i  YG      ]  , , ��  YG ��  ^) �  ^) �  YG ��  YG      ]  , , �  R{ �  W] �?  W] �?  R{ �  R{      ]  , , �-  R{ �-  W] ��  W] ��  R{ �-  R{      ]  , , ��  R{ ��  W]  {  W]  {  R{ ��  R{      ]  , , ��  F� ��  Ki �  Ki �  F� ��  F�      ]  , , �  F� �  Ki �?  Ki �?  F� �  F�      ]  , , �-  F� �-  Ki ��  Ki ��  F� �-  F�      ]  , , ��  F� ��  Ki  {  Ki  {  F� ��  F�      ]  , , i  F� i  Ki   Ki   F� i  F�      ]  , ,   F�   Ki �  Ki �  F�   F�      ]  , , i  R{ i  W]   W]   R{ i  R{      ]  , , ��  R{ ��  W] �  W] �  R{ ��  R{      ]  , , �  R{ �  W] �  W] �  R{ �  R{      ]  , , �  R{ �  W] �S  W] �S  R{ �  R{      ]  , , �A  R{ �A  W] ��  W] ��  R{ �A  R{      ]  , , �{  F� �{  Ki �+  Ki �+  F� �{  F�      ]  , , �  F� �  Ki ��  Ki ��  F� �  F�      ]  , , ��  F� ��  Ki �g  Ki �g  F� ��  F�      ]  , , �U  F� �U  Ki   Ki   F� �U  F�      ]  , , �  F� �  Ki 
�  Ki 
�  F� �  F�      ]  , , �  F� �  Ki A  Ki A  F� �  F�      ]  , ,  �  R{  �  W] �  W] �  R{  �  R{      ]  , , �g  R{ �g  W] �  W] �  R{ �g  R{      ]  , , �  R{ �  W] ��  W] ��  R{ �  R{      ]  , , ��  R{ ��  W] �g  W] �g  R{ ��  R{      ]  , , �U  R{ �U  W]   W]   R{ �U  R{      ]  , , �g  F� �g  Ki �  Ki �  F� �g  F�      ]  , , �  F� �  Ki �  Ki �  F� �  F�      ]  , , �  F� �  Ki �S  Ki �S  F� �  F�      ]  , , �A  F� �A  Ki ��  Ki ��  F� �A  F�      ]  , ,  �  F�  �  Ki �  Ki �  F�  �  F�      ]  , , }  F� }  Ki -  Ki -  F� }  F�      ]  , , �  R{ �  W] 
�  W] 
�  R{ �  R{      ]  , , �{  R{ �{  W] �+  W] �+  R{ �{  R{      ]  , , �  {� �  ~; �3  ~; �3  {� �  {�      ]  , , �9  {� �9  ~; ��  ~; ��  {� �9  {�      ]  , , ��  {� ��  ~; o  ~; o  {� ��  {�      ]  , , ��  � ��  "3 �  "3 �  � ��  �      ]  , , �  � �  "3 �3  "3 �3  � �  �      ]  , , �9  � �9  "3 ��  "3 ��  � �9  �      ]  , , ��  � ��  "3 o  "3 o  � ��  �      ]  , , u  � u  "3 
  "3 
  � u  �      ]  , , 	  � 	  "3 �  "3 �  � 	  �      ]  , , u  {� u  ~; 
  ~; 
  {� u  {�      ]  , , ��  {� ��  ~; �  ~; �  {� ��  {�      ]  , , ��  YG ��  ^) A  ^) A  YG ��  YG      ]  , , �g  ?� �g  D� �  D� �  ?� �g  ?�      ]  , , ��  R{ ��  W] A  W] A  R{ ��  R{      ]  , , ��  F� ��  Ki A  Ki A  F� ��  F�      ]  , , ��  ?� ��  D� A  D� A  ?� ��  ?�      ]  , , �U  YG �U  ^)   ^)   YG �U  YG      ]  , , �  YG �  ^) ��  ^) ��  YG �  YG      ]  , , �  ?� �  D� �  D� �  ?� �  ?�      ]  , , �A  ?� �A  D� ��  D� ��  ?� �A  ?�      ]  , , }  ?� }  D� -  D� -  ?� }  ?�      ]  , , ��  R{ ��  W] �  W] �  R{ ��  R{      ]  , , �{  YG �{  ^) �+  ^) �+  YG �{  YG      ]  , , 
�  YG 
�  ^) �  ^) �  YG 
�  YG      ]  , , �  YG �  ^) �  ^) �  YG �  YG      ]  , , y  YG y  ^) a  ^) a  YG y  YG      ]  , , ;  YG ;  ^) #  ^) #  YG ;  YG      ]  , , �  ?� �  D� �S  D� �S  ?� �  ?�      ]  , , �  YG �  ^) 
�  ^) 
�  YG �  YG      ]  , , ��  YG ��  ^) �g  ^) �g  YG ��  YG      ]  , ,  �  ?�  �  D� �  D� �  ?�  �  ?�      ]  , , �g  ?� �g  D� �  D� �  ?� �g  ?�      @   , ߒ  {z ߒ  ~r �  ~r �  {z ߒ  {z      @   , �,  {z �,  ~r �.  ~r �.  {z �,  {z      @   , 8  o� 8  r P  r P  o� 8  o�      @   , �)  o� �)  {� �A  {� �A  o� �)  o�      @   , �)  c� �)  ~r �S  ~r �S  c� �)  c�      @   , W  c� W  ~r �  ~r �  c� W  c�      @   , �)  r �)  :H �  :H �  r �)  r      @   , �  d� �  o�   o�   d� �  d�      @   , I  d� I  o� �  o� �  d� I  d�      @   , �  d� �  o� �  o� �  d� �  d�      @   , 
  d� 
  o� S  o� S  d� 
  d�      @   , �Q  c� �Q  ~r �}  ~r �}  c� �Q  c�      @   , ��  c� ��  ~r �  ~r �  c� ��  c�      @   , ��  c� ��  ~r �  ~r �  c� ��  c�      @   , �  r �  :H ��  :H ��  r �  r      @   , �Q  r �Q  :H �}  :H �}  r �Q  r      @   , ��  r ��  :H �  :H �  r ��  r      @   , ��  r ��  :H �  :H �  r ��  r      @   ,  +  r  +  :H W  :H W  r  +  r      @   , �  r �  :H �  :H �  r �  r      @   ,  +  c�  +  ~r W  ~r W  c�  +  c�      @   , �  c� �  ~r ��  ~r ��  c� �  c�      @   , �d  {z �d  ~r �j  ~r �j  {z �d  {z      @   , �  {z �  ~r �  ~r �  {z �  {z      @   , ��  {z ��  ~r �  ~r �  {z ��  {z      @   , ��  r ��  "j ��  "j ��  r ��  r      @   , �d  r �d  "j �j  "j �j  r �d  r      @   , �  r �  "j �  "j �  r �  r      @   , ��  r ��  "j �  "j �  r ��  r      @   , >  r >  "j 
D  "j 
D  r >  r      @   , �  r �  "j �  "j �  r �  r      @   , >  {z >  ~r 
D  ~r 
D  {z >  {z      @   , ��  {z ��  ~r ��  ~r ��  {z ��  {z      @   , �Q  o� �Q  {� �i  {� �i  o� �Q  o�      @   , ��  o� ��  {� �  {� �  o� ��  o�      @   , ��  o� ��  {� ��  {� ��  o� ��  o�      @   , ��  "$ ��  .@ ��  .@ ��  "$ ��  "$      @   , �e  "$ �e  .@ �}  .@ �}  "$ �e  "$      @   , �  "$ �  .@ �  .@ �  "$ �  "$      @   , ��  "$ ��  .@ �  .@ �  "$ ��  "$      @   , ?  "$ ?  .@ W  .@ W  "$ ?  "$      @   , �  "$ �  .@ �  .@ �  "$ �  "$      @   ,  +  o�  +  {� C  {� C  o�  +  o�      @   , �  o� �  {� ��  {� ��  o� �  o�      @   , ��  o� ��  {� ��  {� ��  o� ��  o�      @   , �y  o� �y  {� ��  {� ��  o� �y  o�      @   , �  o� �  {� /  {� /  o� �  o�      @   , �=  "$ �=  .@ �U  .@ �U  "$ �=  "$      @   , ��  "$ ��  .@ ��  .@ ��  "$ ��  "$      @   , �y  "$ �y  .@ ��  .@ ��  "$ �y  "$      @   , �  "$ �  .@ /  .@ /  "$ �  "$      @   , �  "$ �  .@ �  .@ �  "$ �  "$      @   , 
S  "$ 
S  .@ k  .@ k  "$ 
S  "$      @   , �  o� �  {� �  {� �  o� �  o�      @   , �=  o� �=  {� �U  {� �U  o� �=  o�      @   , �e  o� �e  {� �}  {� �}  o� �e  o�      @   , �  o� �  {� �  {� �  o� �  o�      @   , ��  o� ��  {� �  {� �  o� ��  o�      @   , �  "$ �  .@ ��  .@ ��  "$ �  "$      @   , �Q  "$ �Q  .@ �i  .@ �i  "$ �Q  "$      @   , ��  "$ ��  .@ �  .@ �  "$ ��  "$      @   , ��  "$ ��  .@ ��  .@ ��  "$ ��  "$      @   ,  +  "$  +  .@ C  .@ C  "$  +  "$      @   , �  "$ �  .@ �  .@ �  "$ �  "$      @   , ?  o� ?  {� W  {� W  o� ?  o�      @   , ��  o� ��  {� ��  {� ��  o� ��  o�      @   , ��  c� ��  o� ��  o� ��  c� ��  c�      @   , �y  c� �y  o� ��  o� ��  c� �y  c�      @   , �  c� �  o� /  o� /  c� �  c�      @   , �=  ., �=  :H �U  :H �U  ., �=  .,      @   , ��  ., ��  :H ��  :H ��  ., ��  .,      @   , �y  ., �y  :H ��  :H ��  ., �y  .,      @   , �  ., �  :H /  :H /  ., �  .,      @   , �  ., �  :H �  :H �  ., �  .,      @   , 
S  ., 
S  :H k  :H k  ., 
S  .,      @   , �  c� �  o� �  o� �  c� �  c�      @   , �=  c� �=  o� �U  o� �U  c� �=  c�      C   , ��  N* ��  O� �z  O� �z  N* ��  N*      C   , �F  N* �F  O� ��  O� ��  N* �F  N*      C   , �  |. �  }� �T  }� �T  |. �  |.      C   , �   & �  !� �T  !� �T   & �   &      C   , �  N* �  O� �  O� �  N* �  N*      C   , �  N* �  O� �T  O� �T  N* �  N*      C   , �T  N* �T  O� �  O� �  N* �T  N*      C   , �z  N* �z  O� �  O� �  N* �z  N*      C   , �  N* �  O� �  O� �  N* �  N*      C   , �  N* �  O� �T  O� �T  N* �  N*      C   , �T  N* �T  O� �  O� �  N* �T  N*      C   , �  N* �  O� 	�  O� 	�  N* �  N*      C   , 	�  N* 	�  O� .  O� .  N* 	�  N*      C   , �  N* �  O� 	�  O� 	�  N* �  N*      C   , �z  N* �z  O� �  O� �  N* �z  N*      C   , �j  z �j  z� ��  z� ��  z �j  z      C   , �j  Q6 �j  Q� ��  Q� ��  Q6 �j  Q6      C   , �j  L �j  L� ��  L� ��  L �j  L      C   , �j  #2 �j  #� ��  #� ��  #2 �j  #2      C   , ��  Z_ ��  ] �3  ] �3  Z_ ��  Z_      C   , '  Z_ '  ] �  ] �  Z_ '  Z_      C   , ��  al ��  b� ��  b� ��  al ��  al      C   , <  al <  b� �  b� �  al <  al      C   , �  S� �  VE ��  VE ��  S� �  S�      C   , �  S� �  VE [  VE [  S� �  S�      C   , ��  S� ��  VE �3  VE �3  S� ��  S�      C   , '  S� '  VE �  VE �  S� '  S�      C   , �~  Q6 �~  Q� ��  Q� ��  Q6 �~  Q6      C   ,   Q6   Q� f  Q� f  Q6   Q6      C   , ��  S� ��  VE �3  VE �3  S� ��  S�      C   , '  S� '  VE �  VE �  S� '  S�      C   , ��  S� ��  VE ��  VE ��  S� ��  S�      C   , �  S� �  VE G  VE G  S� �  S�      C   , ��  Q6 ��  Q� �>  Q� �>  Q6 ��  Q6      C   , �  Q6 �  Q� �  Q� �  Q6 �  Q6      C   , ��  S� ��  VE ��  VE ��  S� ��  S�      C   , �  S� �  VE G  VE G  S� �  S�      C   , 	;  S� 	;  VE 	�  VE 	�  S� 	;  S�      C   , �  S� �  VE ��  VE ��  S� �  S�      C   , �  S� �  VE [  VE [  S� �  S�      C   ,    Q6    Q� R  Q� R  Q6    Q6      C   , �  Q6 �  Q� �  Q� �  Q6 �  Q6      C   , �  f� �  m� �  m� �  f� �  f�      C   , �T  |. �T  }� �  }� �  |. �T  |.      C   , }  f� }  m� '  m� '  f� }  f�      C   , �  |. �  }� 	�  }� 	�  |. �  |.      C   , �  f� �  m� e  m� e  f� �  f�      C   , 7  f� 7  m� �  m� �  f� 7  f�      C   , 7  f� 7  m� �  m� �  f� 7  f�      C   , �  f� �  m� e  m� e  f� �  f�      C   , �  f� �  m� �  m� �  f� �  f�      C   , u  f� u  m�   m�   f� u  f�      C   , �  Z_ �  ] ��  ] ��  Z_ �  Z_      C   , �  Z_ �  ] G  ] G  Z_ �  Z_      C   , �  a� �  b� 7  b� 7  a� �  a�      C   , �  n} �  o� �  o� �  n} �  n}      C   , �  Z_ �  ] ��  ] ��  Z_ �  Z_      C   , ��  q� ��  x} �3  x} �3  q� ��  q�      C   , '  q� '  x} �  x} �  q� '  q�      C   , ��  q� ��  x} ��  x} ��  q� ��  q�      C   , �  q� �  x} G  x} G  q� �  q�      C   , ��  z ��  z� �>  z� �>  z ��  z      C   , �  z �  z� �  z� �  z �  z      C   , �  q� �  x} ��  x} ��  q� �  q�      C   , �  q� �  x} [  x} [  q� �  q�      C   , ��  q� ��  x} �3  x} �3  q� ��  q�      C   , '  q� '  x} �  x} �  q� '  q�      C   , �~  z �~  z� ��  z� ��  z �~  z      C   ,   z   z� f  z� f  z   z      C   , ��  q� ��  x} ��  x} ��  q� ��  q�      C   , �  q� �  x} G  x} G  q� �  q�      C   , 	;  q� 	;  x} 	�  x} 	�  q� 	;  q�      C   , �  q� �  x} ��  x} ��  q� �  q�      C   , �  q� �  x} [  x} [  q� �  q�      C   ,    z    z� R  z� R  z    z      C   , �  z �  z� �  z� �  z �  z      C   , �  f� �  m� ��  m� ��  f� �  f�      C   , �  f� �  m� [  m� [  f� �  f�      C   , ��  f� ��  m� �3  m� �3  f� ��  f�      C   , '  f� '  m� �  m� �  f� '  f�      C   , 7  Z_ 7  ] �  ] �  Z_ 7  Z_      C   , }  Z_ }  ] '  ] '  Z_ }  Z_      C   , �  Z_ �  ] �  ] �  Z_ �  Z_      C   , �  Z_ �  ] e  ] e  Z_ �  Z_      C   , u  Z_ u  ]   ]   Z_ u  Z_      C   , �  Z_ �  ] e  ] e  Z_ �  Z_      C   , 7  Z_ 7  ] �  ] �  Z_ 7  Z_      C   , �  Z_ �  ] �  ] �  Z_ �  Z_      C   , �  Z_ �  ] [  ] [  Z_ �  Z_      C   , 	;  Z_ 	;  ] 	�  ] 	�  Z_ 	;  Z_      C   , ��  Z_ ��  ] ��  ] ��  Z_ ��  Z_      C   , ��  ^t ��  _� \  _� \  ^t ��  ^t      C   , �  p5 �  qW �  qW �  p5 �  p5      C   , �  W& �  XH �  XH �  W& �  W&      C   , �  Z_ �  ] [  ] [  Z_ �  Z_      C   , �z  |. �z  }� �  }� �  |. �z  |.      C   , �M  S� �M  VE ��  VE ��  S� �M  S�      C   , ��  S� ��  VE ��  VE ��  S� ��  S�      C   , �a  Z_ �a  ] �  ] �  Z_ �a  Z_      C   , ��  Z_ ��  ] ��  ] ��  Z_ ��  Z_      C   , �  S� �  VE �Y  VE �Y  S� �  S�      C   , �B  Q6 �B  Q� �  Q� �  Q6 �B  Q6      C   , ��  Q6 ��  Q� �*  Q� �*  Q6 ��  Q6      C   , �u  Z_ �u  ] �  ] �  Z_ �u  Z_      C   , ��  Z_ ��  ] ��  ] ��  Z_ ��  Z_      C   , �  Q6 �  Q� ��  Q� ��  Q6 �  Q6      C   , �M  S� �M  VE ��  VE ��  S� �M  S�      C   , �M  q� �M  x} ��  x} ��  q� �M  q�      C   , ��  q� ��  x} ��  x} ��  q� ��  q�      C   , ��  S� ��  VE ��  VE ��  S� ��  S�      C   , ��  q� ��  x} �E  x} �E  q� ��  q�      C   , �  q� �  x} �Y  x} �Y  q� �  q�      C   , ��  q� ��  x} �m  x} �m  q� ��  q�      C   , �a  q� �a  x} �  x} �  q� �a  q�      C   , �9  Z_ �9  ] ��  ] ��  Z_ �9  Z_      C   , �  S� �  VE �Y  VE �Y  S� �  S�      C   , �%  q� �%  x} ��  x} ��  q� �%  q�      C   , �  z �  z� �  z� �  z �  z      C   , �V  z �V  z� ��  z� ��  z �V  z      C   , ��  S� ��  VE �m  VE �m  S� ��  S�      C   , �a  S� �a  VE �  VE �  S� �a  S�      C   , �  z �  z� �d  z� �d  z �  z      C   , ��  q� ��  x} ��  x} ��  q� ��  q�      C   , �u  q� �u  x} �  x} �  q� �u  q�      C   , �M  Z_ �M  ] ��  ] ��  Z_ �M  Z_      C   , ��  Z_ ��  ] ��  ] ��  Z_ ��  Z_      C   , �9  q� �9  x} ��  x} ��  q� �9  q�      C   , �M  q� �M  x} ��  x} ��  q� �M  q�      C   , ��  q� ��  x} ��  x} ��  q� ��  q�      C   , �%  S� �%  VE ��  VE ��  S� �%  S�      C   , �  Q6 �  Q� �  Q� �  Q6 �  Q6      C   , �  q� �  x} �Y  x} �Y  q� �  q�      C   , �B  z �B  z� �  z� �  z �B  z      C   , ��  z ��  z� �*  z� �*  z ��  z      C   , �V  Q6 �V  Q� ��  Q� ��  Q6 �V  Q6      C   , �%  q� �%  x} ��  x} ��  q� �%  q�      C   , �  z �  z� ��  z� ��  z �  z      C   , �a  q� �a  x} �  x} �  q� �a  q�      C   , �  z �  z� ��  z� ��  z �  z      C   , �  Q6 �  Q� �d  Q� �d  Q6 �  Q6      C   , �a  S� �a  VE �  VE �  S� �a  S�      C   , ��  q� ��  x} �m  x} �m  q� ��  q�      C   , ��  q� ��  x} ��  x} ��  q� ��  q�      C   , �u  q� �u  x} �  x} �  q� �u  q�      C   , �  Z_ �  ] �Y  ] �Y  Z_ �  Z_      C   , �b  al �b  b� �  b� �  al �b  al      C   , �9  q� �9  x} ��  x} ��  q� �9  q�      C   , ��  z ��  z� �  z� �  z ��  z      C   , �F  |. �F  }� ��  }� ��  |. �F  |.      C   , �   al �   b� �J  b� �J  al �   al      C   , ��  S� ��  VE �m  VE �m  S� ��  S�      C   , �.  z �.  z� �x  z� �x  z �.  z      C   , ��  f� ��  m� ��  m� ��  f� ��  f�      C   , �u  f� �u  m� �  m� �  f� �u  f�      C   , ��  S� ��  VE ��  VE ��  S� ��  S�      C   , �u  S� �u  VE �  VE �  S� �u  S�      C   , �9  f� �9  m� ��  m� ��  f� �9  f�      C   , �M  f� �M  m� ��  m� ��  f� �M  f�      C   , ��  f� ��  m� ��  m� ��  f� ��  f�      C   , ��  S� ��  VE �E  VE �E  S� ��  S�      C   , �9  Z_ �9  ] ��  ] ��  Z_ �9  Z_      C   , �  f� �  m� �Y  m� �Y  f� �  f�      C   , �9  S� �9  VE ��  VE ��  S� �9  S�      C   , ��  Q6 ��  Q� �  Q� �  Q6 ��  Q6      C   , ��  |. ��  }� �z  }� �z  |. ��  |.      C   , ��  al ��  b� �  b� �  al ��  al      C   , ��  S� ��  VE ��  VE ��  S� ��  S�      C   , �.  Q6 �.  Q� �x  Q� �x  Q6 �.  Q6      C   , �  |. �  }� �  }� �  |. �  |.      C   , �u  S� �u  VE �  VE �  S� �u  S�      C   , �%  S� �%  VE ��  VE ��  S� �%  S�      C   , �u  Z_ �u  ] �  ] �  Z_ �u  Z_      C   , ��  Z_ ��  ] �m  ] �m  Z_ ��  Z_      C   , �9  S� �9  VE ��  VE ��  S� �9  S�      C   , ��  ^t ��  _� �   _� �   ^t ��  ^t      C   , �<  P� �<  R0 �  R0 �  P� �<  P�      C   , ��  %g ��  ,Q ��  ,Q ��  %g ��  %g      C   , �  ;8 �  <x ��  <x ��  ;8 �  ;8      C   , �"  ;8 �"  <x �l  <x �l  ;8 �"  ;8      C   , �9  G� �9  JQ ��  JQ ��  G� �9  G�      C   , ��  G� ��  JQ �m  JQ �m  G� ��  G�      C   , �a  G� �a  JQ �  JQ �  G� �a  G�      C   , �9  %g �9  ,Q ��  ,Q ��  %g �9  %g      C   , ��  %g ��  ,Q ��  ,Q ��  %g ��  %g      C   , �u  %g �u  ,Q �  ,Q �  %g �u  %g      C   , �z   & �z  !� �  !� �   & �z   &      C   , �   & �  !� �  !� �   & �   &      C   , ��  G� ��  JQ ��  JQ ��  G� ��  G�      C   , �u  G� �u  JQ �  JQ �  G� �u  G�      C   , ��  ;8 ��  <x �
  <x �
  ;8 ��  ;8      C   , �  #2 �  #� ��  #� ��  #2 �  #2      C   , �B  #2 �B  #� �  #� �  #2 �B  #2      C   , ��  #2 ��  #� �*  #� �*  #2 ��  #2      C   , �9  @� �9  C� ��  C� ��  @� �9  @�      C   , ��  @� ��  C� ��  C� ��  @� ��  @�      C   , �.  L �.  L� �x  L� �x  L �.  L      C   , ��  L ��  L� �  L� �  L ��  L      C   , �  >b �  ?p �  ?p �  >b �  >b      C   , �%  %g �%  ,Q ��  ,Q ��  %g �%  %g      C   , ��  %g ��  ,Q �m  ,Q �m  %g ��  %g      C   , �a  %g �a  ,Q �  ,Q �  %g �a  %g      C   , �u  @� �u  C� �  C� �  @� �u  @�      C   , �M  @� �M  C� ��  C� ��  @� �M  @�      C   , �  L �  L� ��  L� ��  L �  L      C   , �B  L �B  L� �  L� �  L �B  L      C   , ��  L ��  L� �*  L� �*  L ��  L      C   , �  %g �  ,Q �Y  ,Q �Y  %g �  %g      C   , �M  %g �M  ,Q ��  ,Q ��  %g �M  %g      C   , ��  %g ��  ,Q ��  ,Q ��  %g ��  %g      C   , �%  G� �%  JQ ��  JQ ��  G� �%  G�      C   , ��  G� ��  JQ �m  JQ �m  G� ��  G�      C   , �a  G� �a  JQ �  JQ �  G� �a  G�      C   , ��  @� ��  C� �m  C� �m  @� ��  @�      C   , �9  %g �9  ,Q ��  ,Q ��  %g �9  %g      C   , �  #2 �  #� �d  #� �d  #2 �  #2      C   , �  #2 �  #� �  #� �  #2 �  #2      C   , �V  #2 �V  #� ��  #� ��  #2 �V  #2      C   , ��  %g ��  ,Q ��  ,Q ��  %g ��  %g      C   , �u  %g �u  ,Q �  ,Q �  %g �u  %g      C   , �  G� �  JQ �Y  JQ �Y  G� �  G�      C   , �M  G� �M  JQ ��  JQ ��  G� �M  G�      C   , ��  G� ��  JQ ��  JQ ��  G� ��  G�      C   , �  0 �  7 �Y  7 �Y  0 �  0      C   , �M  0 �M  7 ��  7 ��  0 �M  0      C   , ��  0 ��  7 ��  7 ��  0 ��  0      C   , �  @� �  C� �Y  C� �Y  @� �  @�      C   , �  G� �  JQ �Y  JQ �Y  G� �  G�      C   , ��  %g ��  ,Q �m  ,Q �m  %g ��  %g      C   , �a  %g �a  ,Q �  ,Q �  %g �a  %g      C   , �M  G� �M  JQ ��  JQ ��  G� �M  G�      C   , �9  0 �9  7 ��  7 ��  0 �9  0      C   , ��  0 ��  7 ��  7 ��  0 ��  0      C   , �u  0 �u  7 �  7 �  0 �u  0      C   , ��  G� ��  JQ ��  JQ ��  G� ��  G�      C   , �9  G� �9  JQ ��  JQ ��  G� �9  G�      C   , ��  G� ��  JQ ��  JQ ��  G� ��  G�      C   , �u  G� �u  JQ �  JQ �  G� �u  G�      C   , �.  #2 �.  #� �x  #� �x  #2 �.  #2      C   , ��  #2 ��  #� �  #� �  #2 ��  #2      C   , �  >b �  ?p �n  ?p �n  >b �  >b      C   , �M  @� �M  C� ��  C� ��  @� �M  @�      C   , ��  @� ��  C� ��  C� ��  @� ��  @�      C   , �  L �  L� �d  L� �d  L �  L      C   , ��  @� ��  C� ��  C� ��  @� ��  @�      C   , �  L �  L� �  L� �  L �  L      C   , �V  L �V  L� ��  L� ��  L �V  L      C   , �a  @� �a  C� �  C� �  @� �a  @�      C   , �  %g �  ,Q �Y  ,Q �Y  %g �  %g      C   , �M  %g �M  ,Q ��  ,Q ��  %g �M  %g      C   , �  @� �  C� �Y  C� �Y  @� �  @�      C   , �%  @� �%  C� ��  C� ��  @� �%  @�      C   , ��  >b ��  ?p �H  ?p �H  >b ��  >b      C   , 
&  >b 
&  ?p �  ?p �  >b 
&  >b      C   , O  G� O  JQ �  JQ �  G� O  G�      C   , �  G� �  JQ ��  JQ ��  G� �  G�      C   , �~  #2 �~  #� ��  #� ��  #2 �~  #2      C   ,   #2   #� f  #� f  #2   #2      C   , �  #2 �  #�   #�   #2 �  #2      C   , �  G� �  JQ [  JQ [  G� �  G�      C   , O  G� O  JQ �  JQ �  G� O  G�      C   , ��  @� ��  C� �3  C� �3  @� ��  @�      C   , ��  @� ��  C� ��  C� ��  @� ��  @�      C   , ��  @� ��  C� �3  C� �3  @� ��  @�      C   , �  %g �  ,Q ��  ,Q ��  %g �  %g      C   , �  %g �  ,Q [  ,Q [  %g �  %g      C   , O  %g O  ,Q �  ,Q �  %g O  %g      C   , ��  %g ��  ,Q ��  ,Q ��  %g ��  %g      C   , �  %g �  ,Q G  ,Q G  %g �  %g      C   , 	;  %g 	;  ,Q 	�  ,Q 	�  %g 	;  %g      C   , ��  G� ��  JQ �3  JQ �3  G� ��  G�      C   , '  G� '  JQ �  JQ �  G� '  G�      C   , �  G� �  JQ o  JQ o  G� �  G�      C   , '  @� '  C� �  C� �  @� '  @�      C   , ��  G� ��  JQ ��  JQ ��  G� ��  G�      C   , �  G� �  JQ G  JQ G  G� �  G�      C   , 	;  G� 	;  JQ 	�  JQ 	�  G� 	;  G�      C   , ��  %g ��  ,Q ��  ,Q ��  %g ��  %g      C   , ��  %g ��  ,Q �3  ,Q �3  %g ��  %g      C   , '  %g '  ,Q �  ,Q �  %g '  %g      C   , �  %g �  ,Q o  ,Q o  %g �  %g      C   , �  %g �  ,Q G  ,Q G  %g �  %g      C   , 	;  %g 	;  ,Q 	�  ,Q 	�  %g 	;  %g      C   , �  %g �  ,Q �  ,Q �  %g �  %g      C   , �  G� �  JQ �  JQ �  G� �  G�      C   , �  @� �  C� o  C� o  @� �  @�      C   , ��  G� ��  JQ �3  JQ �3  G� ��  G�      C   , '  G� '  JQ �  JQ �  G� '  G�      C   , ��  L ��  L� �>  L� �>  L ��  L      C   , ��  #2 ��  #� �>  #� �>  #2 ��  #2      C   , �  #2 �  #� �  #� �  #2 �  #2      C   , 
0  #2 
0  #� z  #� z  #2 
0  #2      C   , �  L �  L� �  L� �  L �  L      C   , 
0  L 
0  L� z  L� z  L 
0  L      C   , �  G� �  JQ o  JQ o  G� �  G�      C   ,    #2    #� R  #� R  #2    #2      C   , �  #2 �  #� �  #� �  #2 �  #2      C   , D  #2 D  #� �  #� �  #2 D  #2      C   , �~  L �~  L� ��  L� ��  L �~  L      C   ,   L   L� f  L� f  L   L      C   , ��  0 ��  7 �3  7 �3  0 ��  0      C   , '  0 '  7 �  7 �  0 '  0      C   , �  0 �  7 o  7 o  0 �  0      C   , �  L �  L�   L�   L �  L      C   , 	;  @� 	;  C� 	�  C� 	�  @� 	;  @�      C   ,    L    L� R  L� R  L    L      C   , �  L �  L� �  L� �  L �  L      C   , D  L D  L� �  L� �  L D  L      C   , �T   & �T  !� �  !� �   & �T   &      C   , ��  %g ��  ,Q �3  ,Q �3  %g ��  %g      C   , '  %g '  ,Q �  ,Q �  %g '  %g      C   , �  0 �  7 ��  7 ��  0 �  0      C   , �  0 �  7 [  7 [  0 �  0      C   , O  0 O  7 �  7 �  0 O  0      C   , �  %g �  ,Q o  ,Q o  %g �  %g      C   , �   & �  !� 	�  !� 	�   & �   &      C   , 	�   & 	�  !� .  !� .   & 	�   &      C   , �  @� �  C� ��  C� ��  @� �  @�      C   , �^  ;8 �^  <x  �  <x  �  ;8 �^  ;8      C   , �  ;8 �  <x F  <x F  ;8 �  ;8      C   , �  ;8 �  <x �  <x �  ;8 �  ;8      C   , �  @� �  C� [  C� [  @� �  @�      C   , O  @� O  C� �  C� �  @� O  @�      C   , �  %g �  ,Q ��  ,Q ��  %g �  %g      C   , �  %g �  ,Q [  ,Q [  %g �  %g      C   , O  %g O  ,Q �  ,Q �  %g O  %g      C   , �  @� �  C� o  C� o  @� �  @�      C   , '  @� '  C� �  C� �  @� '  @�      C   , �  G� �  JQ ��  JQ ��  G� �  G�      C   , ��  G� ��  JQ ��  JQ ��  G� ��  G�      C   , �  G� �  JQ G  JQ G  G� �  G�      C   , �  @� �  C� G  C� G  @� �  @�      C   , 	;  G� 	;  JQ 	�  JQ 	�  G� 	;  G�      C   , �  G� �  JQ [  JQ [  G� �  G�      B  , , �X  N� �X  OG �  OG �  N� �X  N�      B  , , �  N� �  OG �h  OG �h  N� �  N�      B  , , ��  N� ��  OG �  OG �  N� ��  N�      B  , , �  N� �  OG �2  OG �2  N� �  N�      B  , , �&  N� �&  OG ��  OG ��  N� �&  N�      B  , , �  N� �  OG �F  OG �F  N� �  N�      B  , , �:  N� �:  OG ��  OG ��  N� �:  N�      B  , , ��  N� ��  OG ��  OG ��  N� ��  N�      B  , ,  v  N�  v  OG    OG    N�  v  N�      B  , ,   N�   OG �  OG �  N�   N�      B  , , �  N� �  OG \  OG \  N� �  N�      B  , , �  N� �  OG n  OG n  N� �  N�      B  , , �L  N� �L  OG ��  OG ��  N� �L  N�      B  , , �>  N� �>  OG ��  OG ��  N� �>  N�      B  , , ��  N� ��  OG ��  OG ��  N� ��  N�      B  , , �z  N� �z  OG �$  OG �$  N� �z  N�      B  , , �H  N� �H  OG ��  OG ��  N� �H  N�      B  , , ��  N� ��  OG �  OG �  N� ��  N�      B  , , ��  N� ��  OG �.  OG �.  N� ��  N�      B  , , �"  N� �"  OG ��  OG ��  N� �"  N�      B  , , �  N� �  OG j  OG j  N� �  N�      B  , , ^  N� ^  OG   OG   N� ^  N�      B  , ,   N�   OG �  OG �  N�   N�      B  , , �  N� �  OG �J  OG �J  N� �  N�      B  , , �  N� �  OG �<  OG �<  N� �  N�      B  , , �0  N� �0  OG ��  OG ��  N� �0  N�      B  , , ��  N� ��  OG �x  OG �x  N� ��  N�      B  , , ��  N� ��  OG �  OG �  N� ��  N�      B  , , �  N� �  OG �<  OG �<  N� �  N�      B  , , �0  N� �0  OG ��  OG ��  N� �0  N�      B  , , ��  N� ��  OG �x  OG �x  N� ��  N�      B  , , l  N� l  OG   OG   N� l  N�      B  , , 
  N� 
  OG �  OG �  N� 
  N�      B  , , l  N� l  OG   OG   N� l  N�      B  , , ��  N� ��  OG �  OG �  N� ��  N�      B  , , ��  N� ��  OG �  OG �  N� ��  N�      B  , , ��  N� ��  OG �.  OG �.  N� ��  N�      B  , , �"  N� �"  OG ��  OG ��  N� �"  N�      B  , , �  N� �  OG �J  OG �J  N� �  N�      B  , , �>  N� �>  OG ��  OG ��  N� �>  N�      B  , , ��  N� ��  OG ��  OG ��  N� ��  N�      B  , , �z  N� �z  OG �$  OG �$  N� �z  N�      B  , ,   N�   OG �  OG �  N�   N�      B  , , �  N� �  OG `  OG `  N� �  N�      B  , , �  N� �  OG j  OG j  N� �  N�      B  , , �H  N� �H  OG ��  OG ��  N� �H  N�      B  , , �:  N� �:  OG ��  OG ��  N� �:  N�      B  , , ��  N� ��  OG ��  OG ��  N� ��  N�      B  , ,  v  N�  v  OG    OG    N�  v  N�      B  , , �L  N� �L  OG ��  OG ��  N� �L  N�      B  , , ��  N� ��  OG �  OG �  N� ��  N�      B  , , �  N� �  OG �2  OG �2  N� �  N�      B  , , �&  N� �&  OG ��  OG ��  N� �&  N�      B  , , �  N� �  OG n  OG n  N� �  N�      B  , , 
b  N� 
b  OG   OG   N� 
b  N�      B  , ,   N�   OG �  OG �  N�   N�      B  , , �  N� �  OG �F  OG �F  N� �  N�      B  , , �  pq �  q E  q E  pq �  pq      B  , , �  pq �  q �  q �  pq �  pq      B  , , C  pq C  q �  q �  pq C  pq      B  , , �  |� �  }K j  }K j  |� �  |�      B  , ,   |�   }K �  }K �  |�   |�      B  , , +  n� +  oY �  oY �  n� +  n�      B  , ,   n�   oY )  oY )  n�   n�      B  , , �  q� �  r� [  r� [  q� �  q�      B  , , �  sK �  s� [  s� [  sK �  sK      B  , , �  t� �  u] [  u] [  t� �  t�      B  , , �  v �  v� [  v� [  v �  v      B  , , �  w� �  x- [  x- [  w� �  w�      B  , , 	;  q� 	;  r� 	�  r� 	�  q� 	;  q�      B  , , �  q� �  r� [  r� [  q� �  q�      B  , , 	;  sK 	;  s� 	�  s� 	�  sK 	;  sK      B  , , �  sK �  s� [  s� [  sK �  sK      B  , , 	;  t� 	;  u] 	�  u] 	�  t� 	;  t�      B  , , �  t� �  u] [  u] [  t� �  t�      B  , , 	;  v 	;  v� 	�  v� 	�  v 	;  v      B  , , �  v �  v� [  v� [  v �  v      B  , , 	;  w� 	;  x- 	�  x- 	�  w� 	;  w�      B  , , �  w� �  x- [  x- [  w� �  w�      B  , , �  z �  z� �  z� �  z �  z      B  , , �  g/ �  g� [  g� [  g/ �  g/      B  , , �  h� �  iA [  iA [  h� �  h�      B  , , �  i� �  j� [  j� [  i� �  i�      B  , , �  kg �  l [  l [  kg �  kg      B  , , �  l� �  my [  my [  l� �  l�      B  , , �  g/ �  g� �  g� �  g/ �  g/      B  , , }  g/ }  g� '  g� '  g/ }  g/      B  , , �  g/ �  g� e  g� e  g/ �  g/      B  , , 7  g/ 7  g� �  g� �  g/ 7  g/      B  , , �  h� �  iA �  iA �  h� �  h�      B  , , }  h� }  iA '  iA '  h� }  h�      B  , , �  h� �  iA e  iA e  h� �  h�      B  , , 7  h� 7  iA �  iA �  h� 7  h�      B  , , �  i� �  j� �  j� �  i� �  i�      B  , , }  i� }  j� '  j� '  i� }  i�      B  , , �  i� �  j� e  j� e  i� �  i�      B  , , 7  i� 7  j� �  j� �  i� 7  i�      B  , , �  kg �  l �  l �  kg �  kg      B  , , }  kg }  l '  l '  kg }  kg      B  , , �  kg �  l e  l e  kg �  kg      B  , , 7  kg 7  l �  l �  kg 7  kg      B  , , �  l� �  my �  my �  l� �  l�      B  , , }  l� }  my '  my '  l� }  l�      B  , , �  l� �  my e  my e  l� �  l�      B  , , 7  l� 7  my �  my �  l� 7  l�      B  , , 7  g/ 7  g� �  g� �  g/ 7  g/      B  , , �  g/ �  g� e  g� e  g/ �  g/      B  , , �  g/ �  g� �  g� �  g/ �  g/      B  , , u  g/ u  g�   g�   g/ u  g/      B  , , 7  h� 7  iA �  iA �  h� 7  h�      B  , , �  h� �  iA e  iA e  h� �  h�      B  , , �  h� �  iA �  iA �  h� �  h�      B  , , u  h� u  iA   iA   h� u  h�      B  , , 7  i� 7  j� �  j� �  i� 7  i�      B  , , �  i� �  j� e  j� e  i� �  i�      B  , , �  i� �  j� �  j� �  i� �  i�      B  , , u  i� u  j�   j�   i� u  i�      B  , , 7  kg 7  l �  l �  kg 7  kg      B  , , �  kg �  l e  l e  kg �  kg      B  , , �  kg �  l �  l �  kg �  kg      B  , , u  kg u  l   l   kg u  kg      B  , , 7  l� 7  my �  my �  l� 7  l�      B  , , �  l� �  my e  my e  l� �  l�      B  , , �  l� �  my �  my �  l� �  l�      B  , , u  l� u  my   my   l� u  l�      B  , , ��  q� ��  r� �3  r� �3  q� ��  q�      B  , , ��  t� ��  u] ��  u] ��  t� ��  t�      B  , , �  t� �  u] G  u] G  t� �  t�      B  , , '  q� '  r� �  r� �  q� '  q�      B  , , �  t� �  u] ��  u] ��  t� �  t�      B  , , ��  q� ��  r� ��  r� ��  q� ��  q�      B  , , ��  v ��  v� ��  v� ��  v ��  v      B  , , �  v �  v� G  v� G  v �  v      B  , , �  q� �  r� G  r� G  q� �  q�      B  , , �  v �  v� ��  v� ��  v �  v      B  , , ��  sK ��  s� �3  s� �3  sK ��  sK      B  , , ��  w� ��  x- ��  x- ��  w� ��  w�      B  , , �  w� �  x- G  x- G  w� �  w�      B  , , '  sK '  s� �  s� �  sK '  sK      B  , , �  w� �  x- ��  x- ��  w� �  w�      B  , , ��  sK ��  s� ��  s� ��  sK ��  sK      B  , ,  X  z  X  z�   z�   z  X  z      B  , , �  sK �  s� G  s� G  sK �  sK      B  , , �  g/ �  g� ��  g� ��  g/ �  g/      B  , , ��  t� ��  u] �3  u] �3  t� ��  t�      B  , , ��  g/ ��  g� �3  g� �3  g/ ��  g/      B  , , '  g/ '  g� �  g� �  g/ '  g/      B  , , �  h� �  iA ��  iA ��  h� �  h�      B  , , '  t� '  u] �  u] �  t� '  t�      B  , , ��  h� ��  iA �3  iA �3  h� ��  h�      B  , , '  h� '  iA �  iA �  h� '  h�      B  , , �  i� �  j� ��  j� ��  i� �  i�      B  , , ��  t� ��  u] ��  u] ��  t� ��  t�      B  , , ��  i� ��  j� �3  j� �3  i� ��  i�      B  , , '  i� '  j� �  j� �  i� '  i�      B  , , �  kg �  l ��  l ��  kg �  kg      B  , , �  t� �  u] G  u] G  t� �  t�      B  , , ��  kg ��  l �3  l �3  kg ��  kg      B  , , '  kg '  l �  l �  kg '  kg      B  , , �  l� �  my ��  my ��  l� �  l�      B  , , ��  v ��  v� �3  v� �3  v ��  v      B  , , ��  l� ��  my �3  my �3  l� ��  l�      B  , , '  l� '  my �  my �  l� '  l�      B  , , '  v '  v� �  v� �  v '  v      B  , , ��  v ��  v� ��  v� ��  v ��  v      B  , , �  v �  v� G  v� G  v �  v      B  , , ��  w� ��  x- �3  x- �3  w� ��  w�      B  , , '  w� '  x- �  x- �  w� '  w�      B  , , ��  w� ��  x- ��  x- ��  w� ��  w�      B  , , �  w� �  x- G  x- G  w� �  w�      B  , , �D  z �D  z� ��  z� ��  z �D  z      B  , , �  z �  z� �  z� �  z �  z      B  , , �  q� �  r� ��  r� ��  q� �  q�      B  , , ��  |� ��  }K �x  }K �x  |� ��  |�      B  , , ��  q� ��  r� �3  r� �3  q� ��  q�      B  , , '  q� '  r� �  r� �  q� '  q�      B  , , �  sK �  s� ��  s� ��  sK �  sK      B  , , l  |� l  }K   }K   |� l  |�      B  , , ��  sK ��  s� �3  s� �3  sK ��  sK      B  , , '  sK '  s� �  s� �  sK '  sK      B  , , �  t� �  u] ��  u] ��  t� �  t�      B  , , �"  |� �"  }K ��  }K ��  |� �"  |�      B  , , ��  t� ��  u] �3  u] �3  t� ��  t�      B  , , '  t� '  u] �  u] �  t� '  t�      B  , , �  v �  v� ��  v� ��  v �  v      B  , , �&  |� �&  }K ��  }K ��  |� �&  |�      B  , , ��  v ��  v� �3  v� �3  v ��  v      B  , , '  v '  v� �  v� �  v '  v      B  , , �  w� �  x- ��  x- ��  w� �  w�      B  , ,  v  |�  v  }K    }K    |�  v  |�      B  , , ��  w� ��  x- �3  x- �3  w� ��  w�      B  , , '  w� '  x- �  x- �  w� '  w�      B  , , ��  z ��  z� �x  z� �x  z ��  z      B  , , l  z l  z�   z�   z l  z      B  , , ��  q� ��  r� ��  r� ��  q� ��  q�      B  , , �  q� �  r� G  r� G  q� �  q�      B  , , �  |� �  }K n  }K n  |� �  |�      B  , , �  q� �  r� ��  r� ��  q� �  q�      B  , , �z  |� �z  }K �$  }K �$  |� �z  |�      B  , , ��  sK ��  s� ��  s� ��  sK ��  sK      B  , , �  sK �  s� G  s� G  sK �  sK      B  , ,   |�   }K �  }K �  |�   |�      B  , , �  sK �  s� ��  s� ��  sK �  sK      B  , ,  X  ^�  X  _P   _P   ^�  X  ^�      B  , , ��  Q6 ��  Q� �x  Q� �x  Q6 ��  Q6      B  , , l  Q6 l  Q�   Q�   Q6 l  Q6      B  , , ��  S� ��  T� �3  T� �3  S� ��  S�      B  , , '  S� '  T� �  T� �  S� '  S�      B  , , ��  S� ��  T� ��  T� ��  S� ��  S�      B  , , �  S� �  T� G  T� G  S� �  S�      B  , , ��  UK ��  U� �3  U� �3  UK ��  UK      B  , , '  UK '  U� �  U� �  UK '  UK      B  , , ��  UK ��  U� ��  U� ��  UK ��  UK      B  , , �  UK �  U� G  U� G  UK �  UK      B  , , �D  Q6 �D  Q� ��  Q� ��  Q6 �D  Q6      B  , , �  Q6 �  Q� �  Q� �  Q6 �  Q6      B  , , ��  S� ��  T� ��  T� ��  S� ��  S�      B  , , �  S� �  T� G  T� G  S� �  S�      B  , , �  S� �  T� ��  T� ��  S� �  S�      B  , , ��  UK ��  U� ��  U� ��  UK ��  UK      B  , , �  UK �  U� G  U� G  UK �  UK      B  , , �  UK �  U� ��  U� ��  UK �  UK      B  , ,  X  Q6  X  Q�   Q�   Q6  X  Q6      B  , , ��  Z� ��  [Y ��  [Y ��  Z� ��  Z�      B  , , ��  \ ��  \� ��  \� ��  \ ��  \      B  , , �  Z� �  [Y ��  [Y ��  Z� �  Z�      B  , , ��  Z� ��  [Y �3  [Y �3  Z� ��  Z�      B  , , '  Z� '  [Y �  [Y �  Z� '  Z�      B  , , �  \ �  \� ��  \� ��  \ �  \      B  , , ��  \ ��  \� �3  \� �3  \ ��  \      B  , , '  \ '  \� �  \� �  \ '  \      B  , , ��  a� ��  ba ��  ba ��  a� ��  a�      B  , , �  a� �  ba 6  ba 6  a� �  a�      B  , , �  S� �  T� ��  T� ��  S� �  S�      B  , , ��  S� ��  T� �3  T� �3  S� ��  S�      B  , , '  S� '  T� �  T� �  S� '  S�      B  , , �  UK �  U� ��  U� ��  UK �  UK      B  , , ��  UK ��  U� �3  U� �3  UK ��  UK      B  , , �  Z� �  [Y ��  [Y ��  Z� �  Z�      B  , , �  Z� �  [Y G  [Y G  Z� �  Z�      B  , , �  \ �  \� ��  \� ��  \ �  \      B  , , �  \ �  \� G  \� G  \ �  \      B  , , '  UK '  U� �  U� �  UK '  UK      B  , , �  Wb �  X �  X �  Wb �  Wb      B  , , R  Wb R  X �  X �  Wb R  Wb      B  , , �  Wb �  X T  X T  Wb �  Wb      B  , , �  \ �  \� e  \� e  \ �  \      B  , , 7  \ 7  \� �  \� �  \ 7  \      B  , , �  \ �  \� �  \� �  \ �  \      B  , , �  Z� �  [Y [  [Y [  Z� �  Z�      B  , , 	;  Z� 	;  [Y 	�  [Y 	�  Z� 	;  Z�      B  , , �  UK �  U� [  U� [  UK �  UK      B  , , �  \ �  \� [  \� [  \ �  \      B  , , 	;  \ 	;  \� 	�  \� 	�  \ 	;  \      B  , , �  S� �  T� [  T� [  S� �  S�      B  , , �  Q6 �  Q� �  Q� �  Q6 �  Q6      B  , , �  Z� �  [Y [  [Y [  Z� �  Z�      B  , , 	;  UK 	;  U� 	�  U� 	�  UK 	;  UK      B  , , 	;  S� 	;  T� 	�  T� 	�  S� 	;  S�      B  , , 7  Z� 7  [Y �  [Y �  Z� 7  Z�      B  , , �  \ �  \� [  \� [  \ �  \      B  , , }  Z� }  [Y '  [Y '  Z� }  Z�      B  , , �  Z� �  [Y �  [Y �  Z� �  Z�      B  , , �  Z� �  [Y e  [Y e  Z� �  Z�      B  , , 7  \ 7  \� �  \� �  \ 7  \      B  , , =  a� =  ba �  ba �  a� =  a�      B  , , }  \ }  \� '  \� '  \ }  \      B  , , �  S� �  T� [  T� [  S� �  S�      B  , , �  \ �  \� �  \� �  \ �  \      B  , , �  \ �  \� e  \� e  \ �  \      B  , , u  Z� u  [Y   [Y   Z� u  Z�      B  , , �  UK �  U� [  U� [  UK �  UK      B  , , �  Z� �  [Y e  [Y e  Z� �  Z�      B  , , 7  Z� 7  [Y �  [Y �  Z� 7  Z�      B  , , �  Z� �  [Y �  [Y �  Z� �  Z�      B  , , u  \ u  \�   \�   \ u  \      B  , , �  a� �  ba �\  ba �\  a� �  a�      B  , , �u  q� �u  r� �  r� �  q� �u  q�      B  , , �:  |� �:  }K ��  }K ��  |� �:  |�      B  , , �M  q� �M  r� ��  r� ��  q� �M  q�      B  , , ��  q� ��  r� ��  r� ��  q� ��  q�      B  , , ��  |� ��  }K ��  }K ��  |� ��  |�      B  , , ��  sK ��  s� ��  s� ��  sK ��  sK      B  , , �u  sK �u  s� �  s� �  sK �u  sK      B  , , �M  sK �M  s� ��  s� ��  sK �M  sK      B  , , ��  sK ��  s� ��  s� ��  sK ��  sK      B  , , ��  t� ��  u] ��  u] ��  t� ��  t�      B  , , �u  t� �u  u] �  u] �  t� �u  t�      B  , , �M  t� �M  u] ��  u] ��  t� �M  t�      B  , , ��  t� ��  u] ��  u] ��  t� ��  t�      B  , , ��  v ��  v� ��  v� ��  v ��  v      B  , , �u  v �u  v� �  v� �  v �u  v      B  , , �M  v �M  v� ��  v� ��  v �M  v      B  , , ��  v ��  v� ��  v� ��  v ��  v      B  , , ��  w� ��  x- ��  x- ��  w� ��  w�      B  , , �u  w� �u  x- �  x- �  w� �u  w�      B  , , �M  w� �M  x- ��  x- ��  w� �M  w�      B  , , ��  w� ��  x- ��  x- ��  w� ��  w�      B  , , �  z �  z� �<  z� �<  z �  z      B  , , �0  z �0  z� ��  z� ��  z �0  z      B  , , �a  q� �a  r� �  r� �  q� �a  q�      B  , , ��  q� ��  r� ��  r� ��  q� ��  q�      B  , , �u  q� �u  r� �  r� �  q� �u  q�      B  , , �a  sK �a  s� �  s� �  sK �a  sK      B  , , ��  sK ��  s� ��  s� ��  sK ��  sK      B  , , �u  sK �u  s� �  s� �  sK �u  sK      B  , , �a  t� �a  u] �  u] �  t� �a  t�      B  , , ��  t� ��  u] ��  u] ��  t� ��  t�      B  , , �u  t� �u  u] �  u] �  t� �u  t�      B  , , �a  v �a  v� �  v� �  v �a  v      B  , , ��  v ��  v� ��  v� ��  v ��  v      B  , , �u  v �u  v� �  v� �  v �u  v      B  , , ��  q� ��  r� ��  r� ��  q� ��  q�      B  , , �a  w� �a  x- �  x- �  w� �a  w�      B  , , ��  w� ��  x- ��  x- ��  w� ��  w�      B  , , �u  w� �u  x- �  x- �  w� �u  w�      B  , , �  z �  z� ��  z� ��  z �  z      B  , , ��  z ��  z� �d  z� �d  z ��  z      B  , , ��  g/ ��  g� ��  g� ��  g/ ��  g/      B  , , �u  g/ �u  g� �  g� �  g/ �u  g/      B  , , �M  g/ �M  g� ��  g� ��  g/ �M  g/      B  , , ��  g/ ��  g� ��  g� ��  g/ ��  g/      B  , , ��  h� ��  iA ��  iA ��  h� ��  h�      B  , , �u  h� �u  iA �  iA �  h� �u  h�      B  , , �M  h� �M  iA ��  iA ��  h� �M  h�      B  , , ��  h� ��  iA ��  iA ��  h� ��  h�      B  , , ��  i� ��  j� ��  j� ��  i� ��  i�      B  , , �u  i� �u  j� �  j� �  i� �u  i�      B  , , �M  i� �M  j� ��  j� ��  i� �M  i�      B  , , ��  i� ��  j� ��  j� ��  i� ��  i�      B  , , ��  kg ��  l ��  l ��  kg ��  kg      B  , , �u  kg �u  l �  l �  kg �u  kg      B  , , �M  q� �M  r� ��  r� ��  q� �M  q�      B  , , ��  q� ��  r� ��  r� ��  q� ��  q�      B  , , �M  kg �M  l ��  l ��  kg �M  kg      B  , , ��  kg ��  l ��  l ��  kg ��  kg      B  , , ��  l� ��  my ��  my ��  l� ��  l�      B  , , �u  l� �u  my �  my �  l� �u  l�      B  , , �M  l� �M  my ��  my ��  l� �M  l�      B  , , ��  l� ��  my ��  my ��  l� ��  l�      B  , , �a  q� �a  r� �  r� �  q� �a  q�      B  , , �M  sK �M  s� ��  s� ��  sK �M  sK      B  , , ��  sK ��  s� ��  s� ��  sK ��  sK      B  , , �  |� �  }K �2  }K �2  |� �  |�      B  , , �a  sK �a  s� �  s� �  sK �a  sK      B  , , �M  t� �M  u] ��  u] ��  t� �M  t�      B  , , ��  t� ��  u] ��  u] ��  t� ��  t�      B  , , �>  |� �>  }K ��  }K ��  |� �>  |�      B  , , ��  |� ��  }K ��  }K ��  |� ��  |�      B  , , �a  t� �a  u] �  u] �  t� �a  t�      B  , , �M  v �M  v� ��  v� ��  v �M  v      B  , , ��  v ��  v� ��  v� ��  v ��  v      B  , , �  |� �  }K �<  }K �<  |� �  |�      B  , , �a  v �a  v� �  v� �  v �a  v      B  , , �0  |� �0  }K ��  }K ��  |� �0  |�      B  , , �M  w� �M  x- ��  x- ��  w� �M  w�      B  , , ��  w� ��  x- ��  x- ��  w� ��  w�      B  , , �a  w� �a  x- �  x- �  w� �a  w�      B  , , ��  |� ��  }K �  }K �  |� ��  |�      B  , , ��  |� ��  }K �.  }K �.  |� ��  |�      B  , , �  z �  z� �P  z� �P  z �  z      B  , , �X  |� �X  }K �  }K �  |� �X  |�      B  , , �  |� �  }K �h  }K �h  |� �  |�      B  , , ��  v ��  v� �m  v� �m  v ��  v      B  , , �  w� �  x- �Y  x- �Y  w� �  w�      B  , , �  t� �  u] �Y  u] �Y  t� �  t�      B  , , �9  q� �9  r� ��  r� ��  q� �9  q�      B  , , �9  kg �9  l ��  l ��  kg �9  kg      B  , , �9  v �9  v� ��  v� ��  v �9  v      B  , , ��  z ��  z� �  z� �  z ��  z      B  , , �  kg �  l �Y  l �Y  kg �  kg      B  , , ��  w� ��  x- �m  x- �m  w� ��  w�      B  , , �  q� �  r� �Y  r� �Y  q� �  q�      B  , , �  q� �  r� �Y  r� �Y  q� �  q�      B  , , ��  q� ��  r� �m  r� �m  q� ��  q�      B  , , �9  l� �9  my ��  my ��  l� �9  l�      B  , , ��  q� ��  r� �m  r� �m  q� ��  q�      B  , , �9  w� �9  x- ��  x- ��  w� �9  w�      B  , , �9  v �9  v� ��  v� ��  v �9  v      B  , , �  l� �  my �Y  my �Y  l� �  l�      B  , , ��  |� ��  }K �  }K �  |� ��  |�      B  , , �%  q� �%  r� ��  r� ��  q� �%  q�      B  , , �  sK �  s� �Y  s� �Y  sK �  sK      B  , , �~  z �~  z� �(  z� �(  z �~  z      B  , , �9  q� �9  r� ��  r� ��  q� �9  q�      B  , , �  sK �  s� �Y  s� �Y  sK �  sK      B  , , ��  sK ��  s� �m  s� �m  sK ��  sK      B  , , �H  |� �H  }K ��  }K ��  |� �H  |�      B  , , �L  |� �L  }K ��  }K ��  |� �L  |�      B  , , �%  sK �%  s� ��  s� ��  sK �%  sK      B  , , �9  g/ �9  g� ��  g� ��  g/ �9  g/      B  , , ��  sK ��  s� �m  s� �m  sK ��  sK      B  , , �  v �  v� �Y  v� �Y  v �  v      B  , , �  g/ �  g� �Y  g� �Y  g/ �  g/      B  , , �  t� �  u] �Y  u] �Y  t� �  t�      B  , , ��  t� ��  u] �m  u] �m  t� ��  t�      B  , , �j  z �j  z� �  z� �  z �j  z      B  , , �%  t� �%  u] ��  u] ��  t� �%  t�      B  , , �9  sK �9  s� ��  s� ��  sK �9  sK      B  , , �9  h� �9  iA ��  iA ��  h� �9  h�      B  , , �  |� �  }K �J  }K �J  |� �  |�      B  , , �9  t� �9  u] ��  u] ��  t� �9  t�      B  , , �  v �  v� �Y  v� �Y  v �  v      B  , , ��  v ��  v� �m  v� �m  v ��  v      B  , , ��  t� ��  u] �m  u] �m  t� ��  t�      B  , , �  h� �  iA �Y  iA �Y  h� �  h�      B  , , �%  v �%  v� ��  v� ��  v �%  v      B  , , �9  w� �9  x- ��  x- ��  w� �9  w�      B  , , �  |� �  }K �F  }K �F  |� �  |�      B  , , ��  |� ��  }K �  }K �  |� ��  |�      B  , , �  w� �  x- �Y  x- �Y  w� �  w�      B  , , ��  w� ��  x- �m  x- �m  w� ��  w�      B  , , �9  i� �9  j� ��  j� ��  i� �9  i�      B  , , �9  t� �9  u] ��  u] ��  t� �9  t�      B  , , �9  sK �9  s� ��  s� ��  sK �9  sK      B  , , �%  w� �%  x- ��  x- ��  w� �%  w�      B  , , �  z �  z� �  z� �  z �  z      B  , , �  i� �  j� �Y  j� �Y  i� �  i�      B  , , ��  q� ��  r� �E  r� �E  q� ��  q�      B  , , �%  q� �%  r� ��  r� ��  q� �%  q�      B  , , ��  sK ��  s� �E  s� �E  sK ��  sK      B  , , �%  sK �%  s� ��  s� ��  sK �%  sK      B  , , ��  t� ��  u] �E  u] �E  t� ��  t�      B  , , �%  t� �%  u] ��  u] ��  t� �%  t�      B  , , ��  v ��  v� �E  v� �E  v ��  v      B  , , �%  v �%  v� ��  v� ��  v �%  v      B  , , ��  w� ��  x- �E  x- �E  w� ��  w�      B  , , �%  w� �%  x- ��  x- ��  w� �%  w�      B  , , ��  z ��  z� �  z� �  z ��  z      B  , , ��  Q6 ��  Q� �6  Q� �6  Q6 ��  Q6      B  , , �  S� �  T� �Y  T� �Y  S� �  S�      B  , , �9  \ �9  \� ��  \� ��  \ �9  \      B  , , ��  S� ��  T� �m  T� �m  S� ��  S�      B  , , �9  \ �9  \� ��  \� ��  \ �9  \      B  , , �  \ �  \� �Y  \� �Y  \ �  \      B  , , �j  Q6 �j  Q� �  Q� �  Q6 �j  Q6      B  , , �  UK �  U� �Y  U� �Y  UK �  UK      B  , , ��  UK ��  U� �m  U� �m  UK ��  UK      B  , , �~  Q6 �~  Q� �(  Q� �(  Q6 �~  Q6      B  , , �  Z� �  [Y �Y  [Y �Y  Z� �  Z�      B  , , �9  Z� �9  [Y ��  [Y ��  Z� �9  Z�      B  , , �  UK �  U� �Y  U� �Y  UK �  UK      B  , , ��  UK ��  U� �m  U� �m  UK ��  UK      B  , , ��  Q6 ��  Q� �  Q� �  Q6 ��  Q6      B  , , �%  S� �%  T� ��  T� ��  S� �%  S�      B  , , �%  UK �%  U� ��  U� ��  UK �%  UK      B  , , �9  S� �9  T� ��  T� ��  S� �9  S�      B  , , �9  UK �9  U� ��  U� ��  UK �9  UK      B  , , ��  S� ��  T� �m  T� �m  S� ��  S�      B  , , �9  Z� �9  [Y ��  [Y ��  Z� �9  Z�      B  , , ��  S� ��  T� �E  T� �E  S� ��  S�      B  , , ��  Z� ��  [Y �m  [Y �m  Z� ��  Z�      B  , , ��  \ ��  \� �m  \� �m  \ ��  \      B  , , ��  UK ��  U� �E  U� �E  UK ��  UK      B  , , �%  UK �%  U� ��  U� ��  UK �%  UK      B  , , �  Q6 �  Q� �  Q� �  Q6 �  Q6      B  , , �  a� �  ba �  ba �  a� �  a�      B  , , �9  S� �9  T� ��  T� ��  S� �9  S�      B  , , �  S� �  T� �Y  T� �Y  S� �  S�      B  , , �%  S� �%  T� ��  T� ��  S� �%  S�      B  , , �9  UK �9  U� ��  U� ��  UK �9  UK      B  , , �  ^� �  _P ��  _P ��  ^� �  ^�      B  , , �  Q6 �  Q� �<  Q� �<  Q6 �  Q6      B  , , �P  a� �P  ba ��  ba ��  a� �P  a�      B  , , ��  Z� ��  [Y ��  [Y ��  Z� ��  Z�      B  , , �u  S� �u  T� �  T� �  S� �u  S�      B  , , ��  UK ��  U� ��  U� ��  UK ��  UK      B  , , �M  S� �M  T� ��  T� ��  S� �M  S�      B  , , ��  S� ��  T� ��  T� ��  S� ��  S�      B  , , ��  Z� ��  [Y ��  [Y ��  Z� ��  Z�      B  , , ��  UK ��  U� ��  U� ��  UK ��  UK      B  , , ��  \ ��  \� ��  \� ��  \ ��  \      B  , , �a  S� �a  T� �  T� �  S� �a  S�      B  , , ��  S� ��  T� ��  T� ��  S� ��  S�      B  , , ��  UK ��  U� ��  U� ��  UK ��  UK      B  , , �u  \ �u  \� �  \� �  \ �u  \      B  , , �u  UK �u  U� �  U� �  UK �u  UK      B  , , �M  \ �M  \� ��  \� ��  \ �M  \      B  , , �  Q6 �  Q� �P  Q� �P  Q6 �  Q6      B  , , �u  UK �u  U� �  U� �  UK �u  UK      B  , , �u  Z� �u  [Y �  [Y �  Z� �u  Z�      B  , , �u  S� �u  T� �  T� �  S� �u  S�      B  , , ��  Z� ��  [Y ��  [Y ��  Z� ��  Z�      B  , , �M  UK �M  U� ��  U� ��  UK �M  UK      B  , , �a  Z� �a  [Y �  [Y �  Z� �a  Z�      B  , , ��  UK ��  U� ��  U� ��  UK ��  UK      B  , , ��  \ ��  \� ��  \� ��  \ ��  \      B  , , �M  S� �M  T� ��  T� ��  S� �M  S�      B  , , �a  \ �a  \� �  \� �  \ �a  \      B  , , ��  S� ��  T� ��  T� ��  S� ��  S�      B  , , �M  Z� �M  [Y ��  [Y ��  Z� �M  Z�      B  , , �u  Z� �u  [Y �  [Y �  Z� �u  Z�      B  , , �M  UK �M  U� ��  U� ��  UK �M  UK      B  , , �a  S� �a  T� �  T� �  S� �a  S�      B  , , �a  UK �a  U� �  U� �  UK �a  UK      B  , , �u  \ �u  \� �  \� �  \ �u  \      B  , , �  Q6 �  Q� ��  Q� ��  Q6 �  Q6      B  , , ��  Q6 ��  Q� �d  Q� �d  Q6 ��  Q6      B  , , ��  \ ��  \� ��  \� ��  \ ��  \      B  , , �0  Q6 �0  Q� ��  Q� ��  Q6 �0  Q6      B  , , �a  UK �a  U� �  U� �  UK �a  UK      B  , , ��  S� ��  T� ��  T� ��  S� ��  S�      B  , , ��  G� ��  H� ��  H� ��  G� ��  G�      B  , , �u  G� �u  H� �  H� �  G� �u  G�      B  , , �a  IW �a  J �  J �  IW �a  IW      B  , , �r  ;� �r  <- �  <- �  ;� �r  ;�      B  , , �  ;� �  <- ��  <- ��  ;� �  ;�      B  , , �a  A# �a  A� �  A� �  A# �a  A#      B  , , ��  A# ��  A� ��  A� ��  A# ��  A#      B  , , �M  IW �M  J ��  J ��  IW �M  IW      B  , , ��  IW ��  J ��  J ��  IW ��  IW      B  , , �  L �  L� �<  L� �<  L �  L      B  , , �0  L �0  L� ��  L� ��  L �0  L      B  , , �M  B� �M  C5 ��  C5 ��  B� �M  B�      B  , , �a  G� �a  H� �  H� �  G� �a  G�      B  , , �M  IW �M  J ��  J ��  IW �M  IW      B  , , ��  IW ��  J ��  J ��  IW ��  IW      B  , , �M  G� �M  H� ��  H� ��  G� �M  G�      B  , , ��  G� ��  H� ��  H� ��  G� ��  G�      B  , , �u  IW �u  J �  J �  IW �u  IW      B  , , ��  IW ��  J ��  J ��  IW ��  IW      B  , , �M  A# �M  A� ��  A� ��  A# �M  A#      B  , , ��  A# ��  A� ��  A� ��  A# ��  A#      B  , , ��  B� ��  C5 ��  C5 ��  B� ��  B�      B  , , �  L �  L� �P  L� �P  L �  L      B  , , ��  B� ��  C5 ��  C5 ��  B� ��  B�      B  , , �a  IW �a  J �  J �  IW �a  IW      B  , , ��  IW ��  J ��  J ��  IW ��  IW      B  , , �u  IW �u  J �  J �  IW �u  IW      B  , , ��  G� ��  H� ��  H� ��  G� ��  G�      B  , , �u  G� �u  H� �  H� �  G� �u  G�      B  , , ��  A# ��  A� ��  A� ��  A# ��  A#      B  , , �M  B� �M  C5 ��  C5 ��  B� �M  B�      B  , , �u  A# �u  A� �  A� �  A# �u  A#      B  , , �M  A# �M  A� ��  A� ��  A# �M  A#      B  , , �a  G� �a  H� �  H� �  G� �a  G�      B  , , �M  G� �M  H� ��  H� ��  G� �M  G�      B  , , ��  G� ��  H� ��  H� ��  G� ��  G�      B  , , ��  B� ��  C5 ��  C5 ��  B� ��  B�      B  , , �  L �  L� ��  L� ��  L �  L      B  , , ��  L ��  L� �d  L� �d  L ��  L      B  , , �u  B� �u  C5 �  C5 �  B� �u  B�      B  , , �a  B� �a  C5 �  C5 �  B� �a  B�      B  , , �  >� �  ?> �  ?> �  >� �  >�      B  , , �j  >� �j  ?> �  ?> �  >� �j  >�      B  , , �9  IW �9  J ��  J ��  IW �9  IW      B  , , ��  IW ��  J �m  J �m  IW ��  IW      B  , , �  G� �  H� �Y  H� �Y  G� �  G�      B  , , �%  B� �%  C5 ��  C5 ��  B� �%  B�      B  , , �9  G� �9  H� ��  H� ��  G� �9  G�      B  , , �  IW �  J �Y  J �Y  IW �  IW      B  , , �  B� �  C5 �Y  C5 �Y  B� �  B�      B  , , �  A# �  A� �Y  A� �Y  A# �  A#      B  , , �9  A# �9  A� ��  A� ��  A# �9  A#      B  , , �%  IW �%  J ��  J ��  IW �%  IW      B  , , �%  G� �%  H� ��  H� ��  G� �%  G�      B  , , ��  G� ��  H� �m  H� �m  G� ��  G�      B  , , ��  B� ��  C5 �m  C5 �m  B� ��  B�      B  , , ��  ;� ��  <- �~  <- �~  ;� ��  ;�      B  , , ��  A# ��  A� �m  A� �m  A# ��  A#      B  , , �  G� �  H� �Y  H� �Y  G� �  G�      B  , , ��  G� ��  H� �m  H� �m  G� ��  G�      B  , , �  A# �  A� �Y  A� �Y  A# �  A#      B  , , �j  L �j  L� �  L� �  L �j  L      B  , , �  L �  L� �  L� �  L �  L      B  , , �%  A# �%  A� ��  A� ��  A# �%  A#      B  , , �9  B� �9  C5 ��  C5 ��  B� �9  B�      B  , , �  IW �  J �Y  J �Y  IW �  IW      B  , , �~  L �~  L� �(  L� �(  L �~  L      B  , , ��  L ��  L� �  L� �  L ��  L      B  , , ��  IW ��  J �m  J �m  IW ��  IW      B  , , �9  IW �9  J ��  J ��  IW �9  IW      B  , , �  B� �  C5 �Y  C5 �Y  B� �  B�      B  , , �9  G� �9  H� ��  H� ��  G� �9  G�      B  , , �  #2 �  #� �  #� �  #2 �  #2      B  , , �9  ' �9  '� ��  '� ��  ' �9  '      B  , , �  )� �  *� �Y  *� �Y  )� �  )�      B  , , �%  (� �%  )1 ��  )1 ��  (� �%  (�      B  , , �  1� �  2} �Y  2} �Y  1� �  1�      B  , , ��  (� ��  )1 �m  )1 �m  (� ��  (�      B  , , �  (� �  )1 �Y  )1 �Y  (� �  (�      B  , , �H   � �H  !C ��  !C ��   � �H   �      B  , , �9  1� �9  2} ��  2} ��  1� �9  1�      B  , , �  +W �  , �Y  , �Y  +W �  +W      B  , , �  6 �  6� �Y  6� �Y  6 �  6      B  , , �9  (� �9  )1 ��  )1 ��  (� �9  (�      B  , , �  0k �  1 �Y  1 �Y  0k �  0k      B  , , ��  %� ��  &a �m  &a �m  %� ��  %�      B  , , �9  +W �9  , ��  , ��  +W �9  +W      B  , , �9  0k �9  1 ��  1 ��  0k �9  0k      B  , , �%  %� �%  &a ��  &a ��  %� �%  %�      B  , , �  ' �  '� �Y  '� �Y  ' �  '      B  , , ��  %� ��  &a �m  &a �m  %� ��  %�      B  , , �9  6 �9  6� ��  6� ��  6 �9  6      B  , , �%  ' �%  '� ��  '� ��  ' �%  '      B  , , ��   � ��  !C �  !C �   � ��   �      B  , , ��  ' ��  '� �m  '� �m  ' ��  '      B  , , ��  +W ��  , �m  , �m  +W ��  +W      B  , , �9  +W �9  , ��  , ��  +W �9  +W      B  , , �9  ' �9  '� ��  '� ��  ' �9  '      B  , , �  4� �  5M �Y  5M �Y  4� �  4�      B  , , ��  ' ��  '� �m  '� �m  ' ��  '      B  , , �9  %� �9  &a ��  &a ��  %� �9  %�      B  , , �  %� �  &a �Y  &a �Y  %� �  %�      B  , , �  %� �  &a �Y  &a �Y  %� �  %�      B  , , �  (� �  )1 �Y  )1 �Y  (� �  (�      B  , , �9  )� �9  *� ��  *� ��  )� �9  )�      B  , , �   � �  !C �J  !C �J   � �   �      B  , , �9  %� �9  &a ��  &a ��  %� �9  %�      B  , , �~  #2 �~  #� �(  #� �(  #2 �~  #2      B  , , �9  4� �9  5M ��  5M ��  4� �9  4�      B  , , ��  )� ��  *� �m  *� �m  )� ��  )�      B  , , ��  #2 ��  #� �  #� �  #2 ��  #2      B  , , �  )� �  *� �Y  *� �Y  )� �  )�      B  , , �  ' �  '� �Y  '� �Y  ' �  '      B  , , �j  #2 �j  #� �  #� �  #2 �j  #2      B  , , �L   � �L  !C ��  !C ��   � �L   �      B  , , �%  +W �%  , ��  , ��  +W �%  +W      B  , , ��  +W ��  , �m  , �m  +W ��  +W      B  , , ��   � ��  !C �  !C �   � ��   �      B  , , �9  (� �9  )1 ��  )1 ��  (� �9  (�      B  , , �  +W �  , �Y  , �Y  +W �  +W      B  , , �  3; �  3� �Y  3� �Y  3; �  3;      B  , , �   � �  !C �F  !C �F   � �   �      B  , , �9  )� �9  *� ��  *� ��  )� �9  )�      B  , , �9  3; �9  3� ��  3� ��  3; �9  3;      B  , , ��  (� ��  )1 �m  )1 �m  (� ��  (�      B  , , �%  )� �%  *� ��  *� ��  )� �%  )�      B  , , ��  )� ��  *� �m  *� �m  )� ��  )�      B  , , ��  1� ��  2} ��  2} ��  1� ��  1�      B  , , �u  1� �u  2} �  2} �  1� �u  1�      B  , , ��   � ��  !C �  !C �   � ��   �      B  , , ��   � ��  !C �.  !C �.   � ��   �      B  , , �M  %� �M  &a ��  &a ��  %� �M  %�      B  , , ��  %� ��  &a ��  &a ��  %� ��  %�      B  , , ��  ' ��  '� ��  '� ��  ' ��  '      B  , , ��  +W ��  , ��  , ��  +W ��  +W      B  , , �M  0k �M  1 ��  1 ��  0k �M  0k      B  , , ��  0k ��  1 ��  1 ��  0k ��  0k      B  , , ��  (� ��  )1 ��  )1 ��  (� ��  (�      B  , , �u  (� �u  )1 �  )1 �  (� �u  (�      B  , , �u  +W �u  , �  , �  +W �u  +W      B  , , ��  ' ��  '� ��  '� ��  ' ��  '      B  , , ��  +W ��  , ��  , ��  +W ��  +W      B  , , �M  4� �M  5M ��  5M ��  4� �M  4�      B  , , ��  0k ��  1 ��  1 ��  0k ��  0k      B  , , �u  0k �u  1 �  1 �  0k �u  0k      B  , , �u  +W �u  , �  , �  +W �u  +W      B  , , ��  4� ��  5M ��  5M ��  4� ��  4�      B  , , �  #2 �  #� ��  #� ��  #2 �  #2      B  , , �M  ' �M  '� ��  '� ��  ' �M  '      B  , , ��  #2 ��  #� �d  #� �d  #2 ��  #2      B  , , ��  ' ��  '� ��  '� ��  ' ��  '      B  , , �a  (� �a  )1 �  )1 �  (� �a  (�      B  , , �u  ' �u  '� �  '� �  ' �u  '      B  , , �M  (� �M  )1 ��  )1 ��  (� �M  (�      B  , , �   � �  !C �<  !C �<   � �   �      B  , , �  #2 �  #� �P  #� �P  #2 �  #2      B  , , �0   � �0  !C ��  !C ��   � �0   �      B  , , ��  4� ��  5M ��  5M ��  4� ��  4�      B  , , �u  4� �u  5M �  5M �  4� �u  4�      B  , , �a  ' �a  '� �  '� �  ' �a  '      B  , , ��  ' ��  '� ��  '� ��  ' ��  '      B  , , �u  ' �u  '� �  '� �  ' �u  '      B  , , �a  +W �a  , �  , �  +W �a  +W      B  , , �M  )� �M  *� ��  *� ��  )� �M  )�      B  , , ��  )� ��  *� ��  *� ��  )� ��  )�      B  , , ��  (� ��  )1 ��  )1 ��  (� ��  (�      B  , , �a  ' �a  '� �  '� �  ' �a  '      B  , , �a  %� �a  &a �  &a �  %� �a  %�      B  , , �M  %� �M  &a ��  &a ��  %� �M  %�      B  , , ��  %� ��  &a ��  &a ��  %� ��  %�      B  , , �M  3; �M  3� ��  3� ��  3; �M  3;      B  , , ��  3; ��  3� ��  3� ��  3; ��  3;      B  , , ��  )� ��  *� ��  *� ��  )� ��  )�      B  , , �u  )� �u  *� �  *� �  )� �u  )�      B  , , �a  %� �a  &a �  &a �  %� �a  %�      B  , , �:   � �:  !C ��  !C ��   � �:   �      B  , , ��  %� ��  &a ��  &a ��  %� ��  %�      B  , , �u  %� �u  &a �  &a �  %� �u  %�      B  , , �>   � �>  !C ��  !C ��   � �>   �      B  , , ��   � ��  !C ��  !C ��   � ��   �      B  , , ��   � ��  !C ��  !C ��   � ��   �      B  , , ��  %� ��  &a ��  &a ��  %� ��  %�      B  , , ��  )� ��  *� ��  *� ��  )� ��  )�      B  , , �M  6 �M  6� ��  6� ��  6 �M  6      B  , , �  #2 �  #� �<  #� �<  #2 �  #2      B  , , �0  #2 �0  #� ��  #� ��  #2 �0  #2      B  , , �a  )� �a  *� �  *� �  )� �a  )�      B  , , ��  3; ��  3� ��  3� ��  3; ��  3;      B  , , �u  3; �u  3� �  3� �  3; �u  3;      B  , , �u  )� �u  *� �  *� �  )� �u  )�      B  , , ��  6 ��  6� ��  6� ��  6 ��  6      B  , , �M  +W �M  , ��  , ��  +W �M  +W      B  , , ��  +W ��  , ��  , ��  +W ��  +W      B  , , �a  +W �a  , �  , �  +W �a  +W      B  , , �u  %� �u  &a �  &a �  %� �u  %�      B  , , �M  )� �M  *� ��  *� ��  )� �M  )�      B  , , ��  (� ��  )1 ��  )1 ��  (� ��  (�      B  , , �u  (� �u  )1 �  )1 �  (� �u  (�      B  , , �   � �  !C �2  !C �2   � �   �      B  , , �M  1� �M  2} ��  2} ��  1� �M  1�      B  , , �M  +W �M  , ��  , ��  +W �M  +W      B  , , ��  +W ��  , ��  , ��  +W ��  +W      B  , , ��  1� ��  2} ��  2} ��  1� ��  1�      B  , , ��  )� ��  *� ��  *� ��  )� ��  )�      B  , , �M  ' �M  '� ��  '� ��  ' �M  '      B  , , �M  (� �M  )1 ��  )1 ��  (� �M  (�      B  , , ��  (� ��  )1 ��  )1 ��  (� ��  (�      B  , , ��  6 ��  6� ��  6� ��  6 ��  6      B  , , �u  6 �u  6� �  6� �  6 �u  6      B  , , �a  )� �a  *� �  *� �  )� �a  )�      B  , , �a  (� �a  )1 �  )1 �  (� �a  (�      B  , , 
�  >� 
�  ?> *  ?> *  >� 
�  >�      B  , , �  IW �  J o  J o  IW �  IW      B  , , 	;  G� 	;  H� 	�  H� 	�  G� 	;  G�      B  , , �  G� �  H� [  H� [  G� �  G�      B  , , O  G� O  H� �  H� �  G� O  G�      B  , , �  G� �  H� [  H� [  G� �  G�      B  , , O  G� O  H� �  H� �  G� O  G�      B  , , �  A# �  A� o  A� o  A# �  A#      B  , , �  G� �  H� o  H� o  G� �  G�      B  , , �  B� �  C5 [  C5 [  B� �  B�      B  , , O  B� O  C5 �  C5 �  B� O  B�      B  , , 	;  G� 	;  H� 	�  H� 	�  G� 	;  G�      B  , , �  G� �  H� �  H� �  G� �  G�      B  , , 
�  L 
�  L� *  L� *  L 
�  L      B  , , �  IW �  J [  J [  IW �  IW      B  , , 
  L 
  L� �  L� �  L 
  L      B  , , O  IW O  J �  J �  IW O  IW      B  , , L  ;� L  <- �  <- �  ;� L  ;�      B  , , �  ;� �  <- �  <- �  ;� �  ;�      B  , , �  L �  L� �  L� �  L �  L      B  , , �  L �  L� >  L� >  L �  L      B  , , �  IW �  J [  J [  IW �  IW      B  , , �  B� �  C5 o  C5 o  B� �  B�      B  , , 	;  B� 	;  C5 	�  C5 	�  B� 	;  B�      B  , , O  IW O  J �  J �  IW O  IW      B  , , �  A# �  A� o  A� o  A# �  A#      B  , , �  B� �  C5 o  C5 o  B� �  B�      B  , , 	;  A# 	;  A� 	�  A� 	�  A# 	;  A#      B  , , 	;  IW 	;  J 	�  J 	�  IW 	;  IW      B  , , �  G� �  H� o  H� o  G� �  G�      B  , , �  A# �  A� [  A� [  A# �  A#      B  , , O  A# O  A� �  A� �  A# O  A#      B  , , �  IW �  J o  J o  IW �  IW      B  , , 	;  IW 	;  J 	�  J 	�  IW 	;  IW      B  , , �  IW �  J �  J �  IW �  IW      B  , , �D  >� �D  ?> ��  ?> ��  >� �D  >�      B  , , �  G� �  H� G  H� G  G� �  G�      B  , , ��  ;� ��  <-  X  <-  X  ;� ��  ;�      B  , , ��  G� ��  H� �3  H� �3  G� ��  G�      B  , , '  G� '  H� �  H� �  G� '  G�      B  , ,  X  L  X  L�   L�   L  X  L      B  , , '  IW '  J �  J �  IW '  IW      B  , , '  A# '  A� �  A� �  A# '  A#      B  , , �  B� �  C5 G  C5 G  B� �  B�      B  , , '  B� '  C5 �  C5 �  B� '  B�      B  , , ��  B� ��  C5 �3  C5 �3  B� ��  B�      B  , , '  B� '  C5 �  C5 �  B� '  B�      B  , , �  IW �  J ��  J ��  IW �  IW      B  , , �  B� �  C5 ��  C5 ��  B� �  B�      B  , , ��  B� ��  C5 �3  C5 �3  B� ��  B�      B  , , �  A# �  A� G  A� G  A# �  A#      B  , , ��  B� ��  C5 ��  C5 ��  B� ��  B�      B  , , �  IW �  J ��  J ��  IW �  IW      B  , , ��  G� ��  H� ��  H� ��  G� ��  G�      B  , , ��  A# ��  A� �3  A� �3  A# ��  A#      B  , , �  G� �  H� G  H� G  G� �  G�      B  , , �  G� �  H� ��  H� ��  G� �  G�      B  , , ��  IW ��  J ��  J ��  IW ��  IW      B  , , �  IW �  J G  J G  IW �  IW      B  , , ��  A# ��  A� ��  A� ��  A# ��  A#      B  , , �  G� �  H� ��  H� ��  G� �  G�      B  , , �D  L �D  L� ��  L� ��  L �D  L      B  , , ��  G� ��  H� �3  H� �3  G� ��  G�      B  , , '  G� '  H� �  H� �  G� '  G�      B  , , �  L �  L� �  L� �  L �  L      B  , , �  A# �  A� ��  A� ��  A# �  A#      B  , , ��  G� ��  H� ��  H� ��  G� ��  G�      B  , , ��  A# ��  A� �3  A� �3  A# ��  A#      B  , , ��  IW ��  J ��  J ��  IW ��  IW      B  , , �  IW �  J G  J G  IW �  IW      B  , , ��  IW ��  J �3  J �3  IW ��  IW      B  , , '  IW '  J �  J �  IW '  IW      B  , , ��  L ��  L� �x  L� �x  L ��  L      B  , , l  L l  L�   L�   L l  L      B  , , '  A# '  A� �  A� �  A# '  A#      B  , , ��  IW ��  J �3  J �3  IW ��  IW      B  , , '  )� '  *� �  *� �  )� '  )�      B  , , �  (� �  )1 ��  )1 ��  (� �  (�      B  , , ��  ' ��  '� ��  '� ��  ' ��  '      B  , , ��  1� ��  2} �3  2} �3  1� ��  1�      B  , , '  1� '  2} �  2} �  1� '  1�      B  , , �  ' �  '� G  '� G  ' �  '      B  , ,  v   �  v  !C    !C     �  v   �      B  , , ��  #2 ��  #� �x  #� �x  #2 ��  #2      B  , , l  #2 l  #�   #�   #2 l  #2      B  , , �  1� �  2} ��  2} ��  1� �  1�      B  , , ��  ' ��  '� �3  '� �3  ' ��  '      B  , , ��  %� ��  &a �3  &a �3  %� ��  %�      B  , , �  6 �  6� ��  6� ��  6 �  6      B  , , '  %� '  &a �  &a �  %� '  %�      B  , , ��  ' ��  '� �3  '� �3  ' ��  '      B  , , �  %� �  &a ��  &a ��  %� �  %�      B  , , ��  0k ��  1 �3  1 �3  0k ��  0k      B  , , '  0k '  1 �  1 �  0k '  0k      B  , , ��  +W ��  , ��  , ��  +W ��  +W      B  , , �  +W �  , G  , G  +W �  +W      B  , , '  ' '  '� �  '� �  ' '  '      B  , , '  ' '  '� �  '� �  ' '  '      B  , , ��  )� ��  *� ��  *� ��  )� ��  )�      B  , , �"   � �"  !C ��  !C ��   � �"   �      B  , , �  0k �  1 ��  1 ��  0k �  0k      B  , , �  )� �  *� G  *� G  )� �  )�      B  , , ��  +W ��  , �3  , �3  +W ��  +W      B  , , '  +W '  , �  , �  +W '  +W      B  , , ��  (� ��  )1 �3  )1 �3  (� ��  (�      B  , , ��  4� ��  5M �3  5M �3  4� ��  4�      B  , , ��  %� ��  &a ��  &a ��  %� ��  %�      B  , , �  %� �  &a G  &a G  %� �  %�      B  , , '  4� '  5M �  5M �  4� '  4�      B  , , ��  (� ��  )1 ��  )1 ��  (� ��  (�      B  , , �  (� �  )1 G  )1 G  (� �  (�      B  , , �  ' �  '� ��  '� ��  ' �  '      B  , , '  (� '  )1 �  )1 �  (� '  (�      B  , , �  4� �  5M ��  5M ��  4� �  4�      B  , , �D  #2 �D  #� ��  #� ��  #2 �D  #2      B  , , �  #2 �  #� �  #� �  #2 �  #2      B  , , �  )� �  *� ��  *� ��  )� �  )�      B  , , �&   � �&  !C ��  !C ��   � �&   �      B  , , ��  )� ��  *� ��  *� ��  )� ��  )�      B  , , �  )� �  *� G  *� G  )� �  )�      B  , , ��  %� ��  &a ��  &a ��  %� ��  %�      B  , , �  %� �  &a G  &a G  %� �  %�      B  , , �  )� �  *� ��  *� ��  )� �  )�      B  , , ��   � ��  !C �x  !C �x   � ��   �      B  , ,  X  #2  X  #�   #�   #2  X  #2      B  , , l   � l  !C   !C    � l   �      B  , , ��  )� ��  *� �3  *� �3  )� ��  )�      B  , , '  )� '  *� �  *� �  )� '  )�      B  , , ��  %� ��  &a �3  &a �3  %� ��  %�      B  , , ��  3; ��  3� �3  3� �3  3; ��  3;      B  , , '  3; '  3� �  3� �  3; '  3;      B  , , '  %� '  &a �  &a �  %� '  %�      B  , , �  +W �  , ��  , ��  +W �  +W      B  , , ��  +W ��  , �3  , �3  +W ��  +W      B  , , ��  (� ��  )1 ��  )1 ��  (� ��  (�      B  , , �  (� �  )1 G  )1 G  (� �  (�      B  , , '  +W '  , �  , �  +W '  +W      B  , , �  ' �  '� ��  '� ��  ' �  '      B  , , �   � �  !C n  !C n   � �   �      B  , , �  (� �  )1 ��  )1 ��  (� �  (�      B  , , ��  6 ��  6� �3  6� �3  6 ��  6      B  , , �z   � �z  !C �$  !C �$   � �z   �      B  , , ��  (� ��  )1 �3  )1 �3  (� ��  (�      B  , , '  (� '  )1 �  )1 �  (� '  (�      B  , ,    �   !C �  !C �   �    �      B  , , �  +W �  , ��  , ��  +W �  +W      B  , , ��  +W ��  , ��  , ��  +W ��  +W      B  , , �  +W �  , G  , G  +W �  +W      B  , , ��  ' ��  '� ��  '� ��  ' ��  '      B  , , �  ' �  '� G  '� G  ' �  '      B  , , �  3; �  3� ��  3� ��  3; �  3;      B  , , '  6 '  6� �  6� �  6 '  6      B  , , ��  )� ��  *� �3  *� �3  )� ��  )�      B  , , �  %� �  &a ��  &a ��  %� �  %�      B  , , �  (� �  )1 o  )1 o  (� �  (�      B  , , 	;  )� 	;  *� 	�  *� 	�  )� 	;  )�      B  , , �  6 �  6� o  6� o  6 �  6      B  , , �  3; �  3� [  3� [  3; �  3;      B  , , �  +W �  , o  , o  +W �  +W      B  , , O  3; O  3� �  3� �  3; O  3;      B  , , �  4� �  5M o  5M o  4� �  4�      B  , , O  (� O  )1 �  )1 �  (� O  (�      B  , , �  )� �  *� �  *� �  )� �  )�      B  , , 	;  %� 	;  &a 	�  &a 	�  %� 	;  %�      B  , , �  %� �  &a �  &a �  %� �  %�      B  , , �  %� �  &a [  &a [  %� �  %�      B  , , O  %� O  &a �  &a �  %� O  %�      B  , , 	;  (� 	;  )1 	�  )1 	�  (� 	;  (�      B  , , �  (� �  )1 �  )1 �  (� �  (�      B  , , 	;  %� 	;  &a 	�  &a 	�  %� 	;  %�      B  , , �  ' �  '� [  '� [  ' �  '      B  , , O  ' O  '� �  '� �  ' O  '      B  , , �  1� �  2} o  2} o  1� �  1�      B  , , O  )� O  *� �  *� �  )� O  )�      B  , , 	;  ' 	;  '� 	�  '� 	�  ' 	;  '      B  , , 	;  )� 	;  *� 	�  *� 	�  )� 	;  )�      B  , , �  ' �  '� �  '� �  ' �  '      B  , , �  (� �  )1 [  )1 [  (� �  (�      B  , ,    �   !C �  !C �   �    �      B  , , �  4� �  5M [  5M [  4� �  4�      B  , , O  4� O  5M �  5M �  4� O  4�      B  , , �  #2 �  #� �  #� �  #2 �  #2      B  , , �  #2 �  #� >  #� >  #2 �  #2      B  , , 
  #2 
  #� �  #� �  #2 
  #2      B  , , O  (� O  )1 �  )1 �  (� O  (�      B  , , �  1� �  2} [  2} [  1� �  1�      B  , , �  )� �  *� o  *� o  )� �  )�      B  , , 
   � 
  !C �  !C �   � 
   �      B  , , O  1� O  2} �  2} �  1� O  1�      B  , , �   � �  !C \  !C \   � �   �      B  , , 
�  #2 
�  #� *  #� *  #2 
�  #2      B  , , �  )� �  *� [  *� [  )� �  )�      B  , , �  %� �  &a o  &a o  %� �  %�      B  , , �  +W �  , [  , [  +W �  +W      B  , , �  6 �  6� [  6� [  6 �  6      B  , , O  6 O  6� �  6� �  6 O  6      B  , , O  )� O  *� �  *� �  )� O  )�      B  , , 	;  (� 	;  )1 	�  )1 	�  (� 	;  (�      B  , , �  %� �  &a [  &a [  %� �  %�      B  , , �  +W �  , o  , o  +W �  +W      B  , , O  +W O  , �  , �  +W O  +W      B  , , �  ' �  '� o  '� o  ' �  '      B  , , 
b   � 
b  !C   !C    � 
b   �      B  , , �  0k �  1 o  1 o  0k �  0k      B  , , �  ' �  '� o  '� o  ' �  '      B  , , �  3; �  3� o  3� o  3; �  3;      B  , , 	;  +W 	;  , 	�  , 	�  +W 	;  +W      B  , , O  %� O  &a �  &a �  %� O  %�      B  , , �  (� �  )1 o  )1 o  (� �  (�      B  , , �  )� �  *� o  *� o  )� �  )�      B  , , �   � �  !C `  !C `   � �   �      B  , , �  %� �  &a o  &a o  %� �  %�      B  , , �  +W �  , [  , [  +W �  +W      B  , , O  +W O  , �  , �  +W O  +W      B  , , �  )� �  *� [  *� [  )� �  )�      B  , , �  ' �  '� [  '� [  ' �  '      B  , , 	;  +W 	;  , 	�  , 	�  +W 	;  +W      B  , , O  ' O  '� �  '� �  ' O  '      B  , , �  0k �  1 [  1 [  0k �  0k      B  , , 	;  ' 	;  '� 	�  '� 	�  ' 	;  '      B  , , �  +W �  , �  , �  +W �  +W      B  , , O  0k O  1 �  1 �  0k O  0k      B  , , �   � �  !C j  !C j   � �   �      B  , , ^   � ^  !C   !C    � ^   �      B  , , �  (� �  )1 [  )1 [  (� �  (�      C  , , �X  N� �X  OG �  OG �  N� �X  N�      C  , , �  N� �  OG �h  OG �h  N� �  N�      C  , , ��  N� ��  OG �l  OG �l  N� ��  N�      C  , , �`  N� �`  OG �
  OG �
  N� �`  N�      C  , , ��  N� ��  OG ��  OG ��  N� ��  N�      C  , , ��  N� ��  OG �n  OG �n  N� ��  N�      C  , , �b  N� �b  OG �  OG �  N� �b  N�      C  , , �   N� �   OG ��  OG ��  N� �   N�      C  , ,  �  N�  �  OG H  OG H  N�  �  N�      C  , , <  N� <  OG �  OG �  N� <  N�      C  , , �  N� �  OG �  OG �  N� �  N�      C  , , �  N� �  OG F  OG F  N� �  N�      C  , , �$  N� �$  OG ��  OG ��  N� �$  N�      C  , , �*  N� �*  OG ��  OG ��  N� �*  N�      C  , , ��  N� ��  OG �r  OG �r  N� ��  N�      C  , , �f  N� �f  OG �  OG �  N� �f  N�      C  , , �\  N� �\  OG �  OG �  N� �\  N�      C  , , ��  N� ��  OG �  OG �  N� ��  N�      C  , , ��  N� ��  OG �B  OG �B  N� ��  N�      C  , , �6  N� �6  OG ��  OG ��  N� �6  N�      C  , , �  N� �  OG ~  OG ~  N� �  N�      C  , , r  N� r  OG   OG   N� r  N�      C  , ,   N�   OG �  OG �  N�   N�      C  , , �  N� �  OG �6  OG �6  N� �  N�      C  , , �  N� �  OG �<  OG �<  N� �  N�      C  , , �0  N� �0  OG ��  OG ��  N� �0  N�      C  , , ��  N� ��  OG �x  OG �x  N� ��  N�      C  , , ��  N� ��  OG �  OG �  N� ��  N�      C  , , �  N� �  OG �<  OG �<  N� �  N�      C  , , �0  N� �0  OG ��  OG ��  N� �0  N�      C  , , ��  N� ��  OG �x  OG �x  N� ��  N�      C  , , l  N� l  OG   OG   N� l  N�      C  , , 
  N� 
  OG �  OG �  N� 
  N�      C  , , l  N� l  OG   OG   N� l  N�      C  , , ��  N� ��  OG �  OG �  N� ��  N�      C  , , ��  N� ��  OG �  OG �  N� ��  N�      C  , , ��  N� ��  OG �B  OG �B  N� ��  N�      C  , , �6  N� �6  OG ��  OG ��  N� �6  N�      C  , , �  N� �  OG �6  OG �6  N� �  N�      C  , , �*  N� �*  OG ��  OG ��  N� �*  N�      C  , , ��  N� ��  OG �r  OG �r  N� ��  N�      C  , , �f  N� �f  OG �  OG �  N� �f  N�      C  , ,   N�   OG �  OG �  N�   N�      C  , , �  N� �  OG L  OG L  N� �  N�      C  , , �  N� �  OG ~  OG ~  N� �  N�      C  , , �\  N� �\  OG �  OG �  N� �\  N�      C  , , �b  N� �b  OG �  OG �  N� �b  N�      C  , , �   N� �   OG ��  OG ��  N� �   N�      C  , ,  �  N�  �  OG H  OG H  N�  �  N�      C  , , �$  N� �$  OG ��  OG ��  N� �$  N�      C  , , ��  N� ��  OG �l  OG �l  N� ��  N�      C  , , �`  N� �`  OG �
  OG �
  N� �`  N�      C  , , ��  N� ��  OG ��  OG ��  N� ��  N�      C  , , �  N� �  OG F  OG F  N� �  N�      C  , , 
:  N� 
:  OG 
�  OG 
�  N� 
:  N�      C  , , <  N� <  OG �  OG �  N� <  N�      C  , , ��  N� ��  OG �n  OG �n  N� ��  N�      C  , , W  pq W  q   q   pq W  pq      C  , , �  pq �  q 1  q 1  pq �  pq      C  , , �  pq �  q �  q �  pq �  pq      C  , , �  |� �  }K ~  }K ~  |� �  |�      C  , , <  |� <  }K �  }K �  |� <  |�      C  , , �  g/ �  g� �  g� �  g/ �  g/      C  , , }  g/ }  g� '  g� '  g/ }  g/      C  , , �  g/ �  g� e  g� e  g/ �  g/      C  , , 7  g/ 7  g� �  g� �  g/ 7  g/      C  , , �  h� �  iA �  iA �  h� �  h�      C  , , }  h� }  iA '  iA '  h� }  h�      C  , , �  h� �  iA e  iA e  h� �  h�      C  , , 7  h� 7  iA �  iA �  h� 7  h�      C  , , �  i� �  j� �  j� �  i� �  i�      C  , , }  i� }  j� '  j� '  i� }  i�      C  , , �  i� �  j� e  j� e  i� �  i�      C  , , 7  i� 7  j� �  j� �  i� 7  i�      C  , , �  kg �  l �  l �  kg �  kg      C  , , }  kg }  l '  l '  kg }  kg      C  , , �  kg �  l e  l e  kg �  kg      C  , , 7  kg 7  l �  l �  kg 7  kg      C  , , �  l� �  my �  my �  l� �  l�      C  , , }  l� }  my '  my '  l� }  l�      C  , , �  l� �  my e  my e  l� �  l�      C  , , 7  l� 7  my �  my �  l� 7  l�      C  , , 7  g/ 7  g� �  g� �  g/ 7  g/      C  , , �  g/ �  g� e  g� e  g/ �  g/      C  , , �  g/ �  g� �  g� �  g/ �  g/      C  , , u  g/ u  g�   g�   g/ u  g/      C  , , 7  h� 7  iA �  iA �  h� 7  h�      C  , , �  h� �  iA e  iA e  h� �  h�      C  , , �  h� �  iA �  iA �  h� �  h�      C  , , u  h� u  iA   iA   h� u  h�      C  , , 7  i� 7  j� �  j� �  i� 7  i�      C  , , �  i� �  j� e  j� e  i� �  i�      C  , , �  i� �  j� �  j� �  i� �  i�      C  , , u  i� u  j�   j�   i� u  i�      C  , , 7  kg 7  l �  l �  kg 7  kg      C  , , �  kg �  l e  l e  kg �  kg      C  , , �  kg �  l �  l �  kg �  kg      C  , , u  kg u  l   l   kg u  kg      C  , , 7  l� 7  my �  my �  l� 7  l�      C  , , �  l� �  my e  my e  l� �  l�      C  , , �  l� �  my �  my �  l� �  l�      C  , , u  l� u  my   my   l� u  l�      C  , , !  n� !  oY �  oY �  n� !  n�      C  , , �  n� �  oY 3  oY 3  n� �  n�      C  , , �  q� �  r� [  r� [  q� �  q�      C  , , �  sK �  s� [  s� [  sK �  sK      C  , , �  t� �  u] [  u] [  t� �  t�      C  , , �  v �  v� [  v� [  v �  v      C  , , �  w� �  x- [  x- [  w� �  w�      C  , , 	;  q� 	;  r� 	�  r� 	�  q� 	;  q�      C  , , �  q� �  r� [  r� [  q� �  q�      C  , , 	;  sK 	;  s� 	�  s� 	�  sK 	;  sK      C  , , �  sK �  s� [  s� [  sK �  sK      C  , , 	;  t� 	;  u] 	�  u] 	�  t� 	;  t�      C  , , �  t� �  u] [  u] [  t� �  t�      C  , , 	;  v 	;  v� 	�  v� 	�  v 	;  v      C  , , �  v �  v� [  v� [  v �  v      C  , , 	;  w� 	;  x- 	�  x- 	�  w� 	;  w�      C  , , �  w� �  x- [  x- [  w� �  w�      C  , , �  z �  z� �  z� �  z �  z      C  , , �  g/ �  g� [  g� [  g/ �  g/      C  , , �  h� �  iA [  iA [  h� �  h�      C  , , �  i� �  j� [  j� [  i� �  i�      C  , , �  kg �  l [  l [  kg �  kg      C  , , �  l� �  my [  my [  l� �  l�      C  , , '  v '  v� �  v� �  v '  v      C  , , ��  v ��  v� ��  v� ��  v ��  v      C  , , �  v �  v� G  v� G  v �  v      C  , , ��  w� ��  x- �3  x- �3  w� ��  w�      C  , , '  w� '  x- �  x- �  w� '  w�      C  , , ��  w� ��  x- ��  x- ��  w� ��  w�      C  , , �  w� �  x- G  x- G  w� �  w�      C  , , �D  z �D  z� ��  z� ��  z �D  z      C  , , �  z �  z� �  z� �  z �  z      C  , , �  q� �  r� ��  r� ��  q� �  q�      C  , , ��  |� ��  }K �x  }K �x  |� ��  |�      C  , , ��  q� ��  r� �3  r� �3  q� ��  q�      C  , , '  q� '  r� �  r� �  q� '  q�      C  , , �  sK �  s� ��  s� ��  sK �  sK      C  , , l  |� l  }K   }K   |� l  |�      C  , , ��  sK ��  s� �3  s� �3  sK ��  sK      C  , , '  sK '  s� �  s� �  sK '  sK      C  , , �  t� �  u] ��  u] ��  t� �  t�      C  , , �6  |� �6  }K ��  }K ��  |� �6  |�      C  , , ��  t� ��  u] �3  u] �3  t� ��  t�      C  , , '  t� '  u] �  u] �  t� '  t�      C  , , �  v �  v� ��  v� ��  v �  v      C  , , ��  |� ��  }K ��  }K ��  |� ��  |�      C  , , ��  v ��  v� �3  v� �3  v ��  v      C  , , '  v '  v� �  v� �  v '  v      C  , , �  w� �  x- ��  x- ��  w� �  w�      C  , ,  �  |�  �  }K H  }K H  |�  �  |�      C  , , ��  w� ��  x- �3  x- �3  w� ��  w�      C  , , '  w� '  x- �  x- �  w� '  w�      C  , , ��  z ��  z� �x  z� �x  z ��  z      C  , , l  z l  z�   z�   z l  z      C  , , ��  q� ��  r� ��  r� ��  q� ��  q�      C  , , �  q� �  r� G  r� G  q� �  q�      C  , , �  |� �  }K F  }K F  |� �  |�      C  , , �  q� �  r� ��  r� ��  q� �  q�      C  , , �f  |� �f  }K �  }K �  |� �f  |�      C  , , ��  sK ��  s� ��  s� ��  sK ��  sK      C  , , �  sK �  s� G  s� G  sK �  sK      C  , ,   |�   }K �  }K �  |�   |�      C  , , �  sK �  s� ��  s� ��  sK �  sK      C  , , ��  q� ��  r� �3  r� �3  q� ��  q�      C  , , ��  t� ��  u] ��  u] ��  t� ��  t�      C  , , �  t� �  u] G  u] G  t� �  t�      C  , , '  q� '  r� �  r� �  q� '  q�      C  , , �  t� �  u] ��  u] ��  t� �  t�      C  , , ��  q� ��  r� ��  r� ��  q� ��  q�      C  , , ��  v ��  v� ��  v� ��  v ��  v      C  , , �  v �  v� G  v� G  v �  v      C  , , �  q� �  r� G  r� G  q� �  q�      C  , , �  v �  v� ��  v� ��  v �  v      C  , , ��  sK ��  s� �3  s� �3  sK ��  sK      C  , , ��  w� ��  x- ��  x- ��  w� ��  w�      C  , , �  w� �  x- G  x- G  w� �  w�      C  , , '  sK '  s� �  s� �  sK '  sK      C  , , �  w� �  x- ��  x- ��  w� �  w�      C  , , ��  sK ��  s� ��  s� ��  sK ��  sK      C  , ,  X  z  X  z�   z�   z  X  z      C  , , �  sK �  s� G  s� G  sK �  sK      C  , , �  g/ �  g� ��  g� ��  g/ �  g/      C  , , ��  t� ��  u] �3  u] �3  t� ��  t�      C  , , ��  g/ ��  g� �3  g� �3  g/ ��  g/      C  , , '  g/ '  g� �  g� �  g/ '  g/      C  , , �  h� �  iA ��  iA ��  h� �  h�      C  , , '  t� '  u] �  u] �  t� '  t�      C  , , ��  h� ��  iA �3  iA �3  h� ��  h�      C  , , '  h� '  iA �  iA �  h� '  h�      C  , , �  i� �  j� ��  j� ��  i� �  i�      C  , , ��  t� ��  u] ��  u] ��  t� ��  t�      C  , , ��  i� ��  j� �3  j� �3  i� ��  i�      C  , , '  i� '  j� �  j� �  i� '  i�      C  , , �  kg �  l ��  l ��  kg �  kg      C  , , �  t� �  u] G  u] G  t� �  t�      C  , , ��  kg ��  l �3  l �3  kg ��  kg      C  , , '  kg '  l �  l �  kg '  kg      C  , , �  l� �  my ��  my ��  l� �  l�      C  , , ��  v ��  v� �3  v� �3  v ��  v      C  , , ��  l� ��  my �3  my �3  l� ��  l�      C  , , '  l� '  my �  my �  l� '  l�      C  , ,  X  ^�  X  _P   _P   ^�  X  ^�      C  , , �  S� �  T� ��  T� ��  S� �  S�      C  , , ��  UK ��  U� ��  U� ��  UK ��  UK      C  , , �  UK �  U� G  U� G  UK �  UK      C  , , �  UK �  U� ��  U� ��  UK �  UK      C  , ,  X  Q6  X  Q�   Q�   Q6  X  Q6      C  , , ��  Z� ��  [Y ��  [Y ��  Z� ��  Z�      C  , , ��  \ ��  \� ��  \� ��  \ ��  \      C  , , �  Z� �  [Y ��  [Y ��  Z� �  Z�      C  , , ��  Z� ��  [Y �3  [Y �3  Z� ��  Z�      C  , , '  Z� '  [Y �  [Y �  Z� '  Z�      C  , , �  \ �  \� ��  \� ��  \ �  \      C  , , ��  \ ��  \� �3  \� �3  \ ��  \      C  , , '  \ '  \� �  \� �  \ '  \      C  , , ��  a� ��  ba ��  ba ��  a� ��  a�      C  , , �  a� �  ba 6  ba 6  a� �  a�      C  , , �  S� �  T� ��  T� ��  S� �  S�      C  , , ��  S� ��  T� �3  T� �3  S� ��  S�      C  , , '  S� '  T� �  T� �  S� '  S�      C  , , �  UK �  U� ��  U� ��  UK �  UK      C  , , ��  UK ��  U� �3  U� �3  UK ��  UK      C  , , �  Z� �  [Y ��  [Y ��  Z� �  Z�      C  , , �  Z� �  [Y G  [Y G  Z� �  Z�      C  , , �  \ �  \� ��  \� ��  \ �  \      C  , , �  \ �  \� G  \� G  \ �  \      C  , , '  UK '  U� �  U� �  UK '  UK      C  , , ��  Q6 ��  Q� �x  Q� �x  Q6 ��  Q6      C  , , l  Q6 l  Q�   Q�   Q6 l  Q6      C  , , ��  S� ��  T� �3  T� �3  S� ��  S�      C  , , '  S� '  T� �  T� �  S� '  S�      C  , , ��  S� ��  T� ��  T� ��  S� ��  S�      C  , , �  S� �  T� G  T� G  S� �  S�      C  , , ��  UK ��  U� �3  U� �3  UK ��  UK      C  , , '  UK '  U� �  U� �  UK '  UK      C  , , ��  UK ��  U� ��  U� ��  UK ��  UK      C  , , �  UK �  U� G  U� G  UK �  UK      C  , , �D  Q6 �D  Q� ��  Q� ��  Q6 �D  Q6      C  , , �  Q6 �  Q� �  Q� �  Q6 �  Q6      C  , , ��  S� ��  T� ��  T� ��  S� ��  S�      C  , , �  S� �  T� G  T� G  S� �  S�      C  , , �  Wb �  X �  X �  Wb �  Wb      C  , , f  Wb f  X   X   Wb f  Wb      C  , , �  Wb �  X @  X @  Wb �  Wb      C  , , �  Z� �  [Y �  [Y �  Z� �  Z�      C  , , 	;  UK 	;  U� 	�  U� 	�  UK 	;  UK      C  , , u  \ u  \�   \�   \ u  \      C  , , �  UK �  U� [  U� [  UK �  UK      C  , , �  \ �  \� e  \� e  \ �  \      C  , , �  Q6 �  Q� �  Q� �  Q6 �  Q6      C  , , �  \ �  \� [  \� [  \ �  \      C  , , 7  \ 7  \� �  \� �  \ 7  \      C  , , �  \ �  \� �  \� �  \ �  \      C  , , �  Z� �  [Y [  [Y [  Z� �  Z�      C  , , 	;  Z� 	;  [Y 	�  [Y 	�  Z� 	;  Z�      C  , , u  Z� u  [Y   [Y   Z� u  Z�      C  , , �  S� �  T� [  T� [  S� �  S�      C  , , �  \ �  \� [  \� [  \ �  \      C  , , 	;  \ 	;  \� 	�  \� 	�  \ 	;  \      C  , , �  Z� �  [Y e  [Y e  Z� �  Z�      C  , , �  UK �  U� [  U� [  UK �  UK      C  , , 	;  S� 	;  T� 	�  T� 	�  S� 	;  S�      C  , , =  a� =  ba �  ba �  a� =  a�      C  , , 7  Z� 7  [Y �  [Y �  Z� 7  Z�      C  , , �  S� �  T� [  T� [  S� �  S�      C  , , 7  Z� 7  [Y �  [Y �  Z� 7  Z�      C  , , }  Z� }  [Y '  [Y '  Z� }  Z�      C  , , �  Z� �  [Y �  [Y �  Z� �  Z�      C  , , �  Z� �  [Y e  [Y e  Z� �  Z�      C  , , 7  \ 7  \� �  \� �  \ 7  \      C  , , }  \ }  \� '  \� '  \ }  \      C  , , �  \ �  \� �  \� �  \ �  \      C  , , �  \ �  \� e  \� e  \ �  \      C  , , �  Z� �  [Y [  [Y [  Z� �  Z�      C  , , �*  |� �*  }K ��  }K ��  |� �*  |�      C  , , �  a� �  ba �\  ba �\  a� �  a�      C  , , �a  sK �a  s� �  s� �  sK �a  sK      C  , , �M  t� �M  u] ��  u] ��  t� �M  t�      C  , , ��  t� ��  u] ��  u] ��  t� ��  t�      C  , , �  |� �  }K �<  }K �<  |� �  |�      C  , , �a  t� �a  u] �  u] �  t� �a  t�      C  , , �0  |� �0  }K ��  }K ��  |� �0  |�      C  , , �M  v �M  v� ��  v� ��  v �M  v      C  , , ��  v ��  v� ��  v� ��  v ��  v      C  , , �a  v �a  v� �  v� �  v �a  v      C  , , ��  |� ��  }K �  }K �  |� ��  |�      C  , , ��  |� ��  }K �B  }K �B  |� ��  |�      C  , , �M  w� �M  x- ��  x- ��  w� �M  w�      C  , , ��  w� ��  x- ��  x- ��  w� ��  w�      C  , , �a  w� �a  x- �  x- �  w� �a  w�      C  , , �b  |� �b  }K �  }K �  |� �b  |�      C  , , �  z �  z� �P  z� �P  z �  z      C  , , �   |� �   }K ��  }K ��  |� �   |�      C  , , ��  q� ��  r� ��  r� ��  q� ��  q�      C  , , �u  q� �u  r� �  r� �  q� �u  q�      C  , , �M  q� �M  r� ��  r� ��  q� �M  q�      C  , , ��  q� ��  r� ��  r� ��  q� ��  q�      C  , , ��  sK ��  s� ��  s� ��  sK ��  sK      C  , , �u  sK �u  s� �  s� �  sK �u  sK      C  , , �M  sK �M  s� ��  s� ��  sK �M  sK      C  , , ��  sK ��  s� ��  s� ��  sK ��  sK      C  , , ��  t� ��  u] ��  u] ��  t� ��  t�      C  , , �u  t� �u  u] �  u] �  t� �u  t�      C  , , �M  t� �M  u] ��  u] ��  t� �M  t�      C  , , ��  t� ��  u] ��  u] ��  t� ��  t�      C  , , ��  v ��  v� ��  v� ��  v ��  v      C  , , �u  v �u  v� �  v� �  v �u  v      C  , , �M  v �M  v� ��  v� ��  v �M  v      C  , , ��  v ��  v� ��  v� ��  v ��  v      C  , , ��  w� ��  x- ��  x- ��  w� ��  w�      C  , , �u  w� �u  x- �  x- �  w� �u  w�      C  , , �M  w� �M  x- ��  x- ��  w� �M  w�      C  , , ��  w� ��  x- ��  x- ��  w� ��  w�      C  , , �  z �  z� �<  z� �<  z �  z      C  , , �0  z �0  z� ��  z� ��  z �0  z      C  , , �a  q� �a  r� �  r� �  q� �a  q�      C  , , ��  |� ��  }K �r  }K �r  |� ��  |�      C  , , ��  q� ��  r� ��  r� ��  q� ��  q�      C  , , �u  q� �u  r� �  r� �  q� �u  q�      C  , , �a  sK �a  s� �  s� �  sK �a  sK      C  , , ��  sK ��  s� ��  s� ��  sK ��  sK      C  , , �u  sK �u  s� �  s� �  sK �u  sK      C  , , �a  t� �a  u] �  u] �  t� �a  t�      C  , , ��  t� ��  u] ��  u] ��  t� ��  t�      C  , , �u  t� �u  u] �  u] �  t� �u  t�      C  , , �a  v �a  v� �  v� �  v �a  v      C  , , ��  v ��  v� ��  v� ��  v ��  v      C  , , �u  v �u  v� �  v� �  v �u  v      C  , , �a  w� �a  x- �  x- �  w� �a  w�      C  , , ��  w� ��  x- ��  x- ��  w� ��  w�      C  , , �u  w� �u  x- �  x- �  w� �u  w�      C  , , �  z �  z� ��  z� ��  z �  z      C  , , ��  z ��  z� �d  z� �d  z ��  z      C  , , ��  g/ ��  g� ��  g� ��  g/ ��  g/      C  , , �u  g/ �u  g� �  g� �  g/ �u  g/      C  , , �M  g/ �M  g� ��  g� ��  g/ �M  g/      C  , , ��  g/ ��  g� ��  g� ��  g/ ��  g/      C  , , ��  h� ��  iA ��  iA ��  h� ��  h�      C  , , �u  h� �u  iA �  iA �  h� �u  h�      C  , , �M  h� �M  iA ��  iA ��  h� �M  h�      C  , , ��  h� ��  iA ��  iA ��  h� ��  h�      C  , , ��  i� ��  j� ��  j� ��  i� ��  i�      C  , , �u  i� �u  j� �  j� �  i� �u  i�      C  , , �M  q� �M  r� ��  r� ��  q� �M  q�      C  , , ��  q� ��  r� ��  r� ��  q� ��  q�      C  , , �M  i� �M  j� ��  j� ��  i� �M  i�      C  , , ��  i� ��  j� ��  j� ��  i� ��  i�      C  , , �`  |� �`  }K �
  }K �
  |� �`  |�      C  , , ��  kg ��  l ��  l ��  kg ��  kg      C  , , �u  kg �u  l �  l �  kg �u  kg      C  , , �M  kg �M  l ��  l ��  kg �M  kg      C  , , ��  kg ��  l ��  l ��  kg ��  kg      C  , , �a  q� �a  r� �  r� �  q� �a  q�      C  , , ��  l� ��  my ��  my ��  l� ��  l�      C  , , �u  l� �u  my �  my �  l� �u  l�      C  , , �M  l� �M  my ��  my ��  l� �M  l�      C  , , ��  l� ��  my ��  my ��  l� ��  l�      C  , , �M  sK �M  s� ��  s� ��  sK �M  sK      C  , , ��  sK ��  s� ��  s� ��  sK ��  sK      C  , , �  |� �  }K �h  }K �h  |� �  |�      C  , , �X  |� �X  }K �  }K �  |� �X  |�      C  , , �9  t� �9  u] ��  u] ��  t� �9  t�      C  , , �9  t� �9  u] ��  u] ��  t� �9  t�      C  , , ��  v ��  v� �m  v� �m  v ��  v      C  , , �\  |� �\  }K �  }K �  |� �\  |�      C  , , �%  sK �%  s� ��  s� ��  sK �%  sK      C  , , �9  v �9  v� ��  v� ��  v �9  v      C  , , �  t� �  u] �Y  u] �Y  t� �  t�      C  , , ��  w� ��  x- �m  x- �m  w� ��  w�      C  , , �%  w� �%  x- ��  x- ��  w� �%  w�      C  , , �  z �  z� �  z� �  z �  z      C  , , �9  w� �9  x- ��  x- ��  w� �9  w�      C  , , �9  v �9  v� ��  v� ��  v �9  v      C  , , ��  |� ��  }K �  }K �  |� ��  |�      C  , , �~  z �~  z� �(  z� �(  z �~  z      C  , , �  v �  v� �Y  v� �Y  v �  v      C  , , �  v �  v� �Y  v� �Y  v �  v      C  , , �9  g/ �9  g� ��  g� ��  g/ �9  g/      C  , , �j  z �j  z� �  z� �  z �j  z      C  , , ��  v ��  v� �m  v� �m  v ��  v      C  , , �  g/ �  g� �Y  g� �Y  g/ �  g/      C  , , �9  w� �9  x- ��  x- ��  w� �9  w�      C  , , �  t� �  u] �Y  u] �Y  t� �  t�      C  , , �9  h� �9  iA ��  iA ��  h� �9  h�      C  , , ��  |� ��  }K �n  }K �n  |� ��  |�      C  , , �  w� �  x- �Y  x- �Y  w� �  w�      C  , , ��  |� ��  }K �l  }K �l  |� ��  |�      C  , , �  h� �  iA �Y  iA �Y  h� �  h�      C  , , �9  q� �9  r� ��  r� ��  q� �9  q�      C  , , ��  t� ��  u] �m  u] �m  t� ��  t�      C  , , ��  z ��  z� �  z� �  z ��  z      C  , , ��  sK ��  s� �m  s� �m  sK ��  sK      C  , , �9  i� �9  j� ��  j� ��  i� �9  i�      C  , , �  q� �  r� �Y  r� �Y  q� �  q�      C  , , ��  q� ��  r� �m  r� �m  q� ��  q�      C  , , �%  v �%  v� ��  v� ��  v �%  v      C  , , �  i� �  j� �Y  j� �Y  i� �  i�      C  , , �  sK �  s� �Y  s� �Y  sK �  sK      C  , , �9  q� �9  r� ��  r� ��  q� �9  q�      C  , , �  q� �  r� �Y  r� �Y  q� �  q�      C  , , ��  q� ��  r� �m  r� �m  q� ��  q�      C  , , �9  kg �9  l ��  l ��  kg �9  kg      C  , , �9  sK �9  s� ��  s� ��  sK �9  sK      C  , , ��  sK ��  s� �m  s� �m  sK ��  sK      C  , , �%  t� �%  u] ��  u] ��  t� �%  t�      C  , , �  kg �  l �Y  l �Y  kg �  kg      C  , , �  w� �  x- �Y  x- �Y  w� �  w�      C  , , �9  sK �9  s� ��  s� ��  sK �9  sK      C  , , �$  |� �$  }K ��  }K ��  |� �$  |�      C  , , �%  q� �%  r� ��  r� ��  q� �%  q�      C  , , �9  l� �9  my ��  my ��  l� �9  l�      C  , , �  sK �  s� �Y  s� �Y  sK �  sK      C  , , ��  t� ��  u] �m  u] �m  t� ��  t�      C  , , ��  w� ��  x- �m  x- �m  w� ��  w�      C  , , �  |� �  }K �6  }K �6  |� �  |�      C  , , �  l� �  my �Y  my �Y  l� �  l�      C  , , ��  q� ��  r� �E  r� �E  q� ��  q�      C  , , �%  q� �%  r� ��  r� ��  q� �%  q�      C  , , ��  sK ��  s� �E  s� �E  sK ��  sK      C  , , �%  sK �%  s� ��  s� ��  sK �%  sK      C  , , ��  t� ��  u] �E  u] �E  t� ��  t�      C  , , �%  t� �%  u] ��  u] ��  t� �%  t�      C  , , ��  v ��  v� �E  v� �E  v ��  v      C  , , �%  v �%  v� ��  v� ��  v �%  v      C  , , ��  w� ��  x- �E  x- �E  w� ��  w�      C  , , �%  w� �%  x- ��  x- ��  w� �%  w�      C  , , ��  z ��  z� �  z� �  z ��  z      C  , , ��  Q6 ��  Q� �6  Q� �6  Q6 ��  Q6      C  , , �  S� �  T� �Y  T� �Y  S� �  S�      C  , , �9  S� �9  T� ��  T� ��  S� �9  S�      C  , , ��  S� ��  T� �m  T� �m  S� ��  S�      C  , , �  UK �  U� �Y  U� �Y  UK �  UK      C  , , �~  Q6 �~  Q� �(  Q� �(  Q6 �~  Q6      C  , , �9  S� �9  T� ��  T� ��  S� �9  S�      C  , , ��  UK ��  U� �m  U� �m  UK ��  UK      C  , , �j  Q6 �j  Q� �  Q� �  Q6 �j  Q6      C  , , �  UK �  U� �Y  U� �Y  UK �  UK      C  , , ��  UK ��  U� �m  U� �m  UK ��  UK      C  , , �9  \ �9  \� ��  \� ��  \ �9  \      C  , , �  a� �  ba �  ba �  a� �  a�      C  , , ��  S� ��  T� �E  T� �E  S� ��  S�      C  , , �9  Z� �9  [Y ��  [Y ��  Z� �9  Z�      C  , , �%  S� �%  T� ��  T� ��  S� �%  S�      C  , , ��  Z� ��  [Y �m  [Y �m  Z� ��  Z�      C  , , ��  UK ��  U� �E  U� �E  UK ��  UK      C  , , �9  \ �9  \� ��  \� ��  \ �9  \      C  , , �%  UK �%  U� ��  U� ��  UK �%  UK      C  , , ��  \ ��  \� �m  \� �m  \ ��  \      C  , , �  Z� �  [Y �Y  [Y �Y  Z� �  Z�      C  , , ��  Q6 ��  Q� �  Q� �  Q6 ��  Q6      C  , , �9  UK �9  U� ��  U� ��  UK �9  UK      C  , , ��  S� ��  T� �m  T� �m  S� ��  S�      C  , , �9  UK �9  U� ��  U� ��  UK �9  UK      C  , , �  \ �  \� �Y  \� �Y  \ �  \      C  , , �%  UK �%  U� ��  U� ��  UK �%  UK      C  , , �9  Z� �9  [Y ��  [Y ��  Z� �9  Z�      C  , , �  Q6 �  Q� �  Q� �  Q6 �  Q6      C  , , �  S� �  T� �Y  T� �Y  S� �  S�      C  , , �%  S� �%  T� ��  T� ��  S� �%  S�      C  , , �  ^� �  _P ��  _P ��  ^� �  ^�      C  , , �u  Z� �u  [Y �  [Y �  Z� �u  Z�      C  , , �M  UK �M  U� ��  U� ��  UK �M  UK      C  , , �a  S� �a  T� �  T� �  S� �a  S�      C  , , ��  UK ��  U� ��  U� ��  UK ��  UK      C  , , ��  \ ��  \� ��  \� ��  \ ��  \      C  , , �a  S� �a  T� �  T� �  S� �a  S�      C  , , ��  \ ��  \� ��  \� ��  \ ��  \      C  , , �u  UK �u  U� �  U� �  UK �u  UK      C  , , ��  Z� ��  [Y ��  [Y ��  Z� ��  Z�      C  , , �u  \ �u  \� �  \� �  \ �u  \      C  , , �u  Z� �u  [Y �  [Y �  Z� �u  Z�      C  , , �M  \ �M  \� ��  \� ��  \ �M  \      C  , , ��  S� ��  T� ��  T� ��  S� ��  S�      C  , , �a  Z� �a  [Y �  [Y �  Z� �a  Z�      C  , , �u  S� �u  T� �  T� �  S� �u  S�      C  , , ��  Z� ��  [Y ��  [Y ��  Z� ��  Z�      C  , , �u  \ �u  \� �  \� �  \ �u  \      C  , , �a  UK �a  U� �  U� �  UK �a  UK      C  , , �  Q6 �  Q� ��  Q� ��  Q6 �  Q6      C  , , ��  Q6 ��  Q� �d  Q� �d  Q6 ��  Q6      C  , , ��  UK ��  U� ��  U� ��  UK ��  UK      C  , , ��  S� ��  T� ��  T� ��  S� ��  S�      C  , , �P  a� �P  ba ��  ba ��  a� �P  a�      C  , , �0  Q6 �0  Q� ��  Q� ��  Q6 �0  Q6      C  , , ��  UK ��  U� ��  U� ��  UK ��  UK      C  , , �u  S� �u  T� �  T� �  S� �u  S�      C  , , �a  \ �a  \� �  \� �  \ �a  \      C  , , �M  Z� �M  [Y ��  [Y ��  Z� �M  Z�      C  , , �M  UK �M  U� ��  U� ��  UK �M  UK      C  , , ��  UK ��  U� ��  U� ��  UK ��  UK      C  , , �M  S� �M  T� ��  T� ��  S� �M  S�      C  , , ��  S� ��  T� ��  T� ��  S� ��  S�      C  , , �a  UK �a  U� �  U� �  UK �a  UK      C  , , �  Q6 �  Q� �<  Q� �<  Q6 �  Q6      C  , , �  Q6 �  Q� �P  Q� �P  Q6 �  Q6      C  , , ��  Z� ��  [Y ��  [Y ��  Z� ��  Z�      C  , , �M  S� �M  T� ��  T� ��  S� �M  S�      C  , , ��  S� ��  T� ��  T� ��  S� ��  S�      C  , , ��  \ ��  \� ��  \� ��  \ ��  \      C  , , �u  UK �u  U� �  U� �  UK �u  UK      C  , , �*   � �*  !C ��  !C ��   � �*   �      C  , , ��  IW ��  J ��  J ��  IW ��  IW      C  , , �u  IW �u  J �  J �  IW �u  IW      C  , , ��  A# ��  A� ��  A� ��  A# ��  A#      C  , , �u  G� �u  H� �  H� �  G� �u  G�      C  , , �a  G� �a  H� �  H� �  G� �a  G�      C  , , �M  A# �M  A� ��  A� ��  A# �M  A#      C  , , �M  B� �M  C5 ��  C5 ��  B� �M  B�      C  , , �M  G� �M  H� ��  H� ��  G� �M  G�      C  , , �  L �  L� ��  L� ��  L �  L      C  , , ��  L ��  L� �d  L� �d  L ��  L      C  , , ��  G� ��  H� ��  H� ��  G� ��  G�      C  , , ��  B� ��  C5 ��  C5 ��  B� ��  B�      C  , , ��  A# ��  A� ��  A� ��  A# ��  A#      C  , , �u  A# �u  A� �  A� �  A# �u  A#      C  , , �a  IW �a  J �  J �  IW �a  IW      C  , , �a  B� �a  C5 �  C5 �  B� �a  B�      C  , , ��  G� ��  H� ��  H� ��  G� ��  G�      C  , , �u  G� �u  H� �  H� �  G� �u  G�      C  , , �M  IW �M  J ��  J ��  IW �M  IW      C  , , ��  IW ��  J ��  J ��  IW ��  IW      C  , , ��  A# ��  A� ��  A� ��  A# ��  A#      C  , , �a  G� �a  H� �  H� �  G� �a  G�      C  , , �  L �  L� �<  L� �<  L �  L      C  , , �0  L �0  L� ��  L� ��  L �0  L      C  , , �r  ;� �r  <- �  <- �  ;� �r  ;�      C  , , �  ;� �  <- ��  <- ��  ;� �  ;�      C  , , �M  G� �M  H� ��  H� ��  G� �M  G�      C  , , ��  G� ��  H� ��  H� ��  G� ��  G�      C  , , ��  B� ��  C5 ��  C5 ��  B� ��  B�      C  , , �u  B� �u  C5 �  C5 �  B� �u  B�      C  , , ��  IW ��  J ��  J ��  IW ��  IW      C  , , �u  IW �u  J �  J �  IW �u  IW      C  , , �  L �  L� �P  L� �P  L �  L      C  , , �a  A# �a  A� �  A� �  A# �a  A#      C  , , �M  IW �M  J ��  J ��  IW �M  IW      C  , , ��  IW ��  J ��  J ��  IW ��  IW      C  , , �a  IW �a  J �  J �  IW �a  IW      C  , , �M  B� �M  C5 ��  C5 ��  B� �M  B�      C  , , ��  B� ��  C5 ��  C5 ��  B� ��  B�      C  , , �M  A# �M  A� ��  A� ��  A# �M  A#      C  , , ��  G� ��  H� ��  H� ��  G� ��  G�      C  , , �  >� �  ?> �  ?> �  >� �  >�      C  , , �j  >� �j  ?> �  ?> �  >� �j  >�      C  , , �9  IW �9  J ��  J ��  IW �9  IW      C  , , �  B� �  C5 �Y  C5 �Y  B� �  B�      C  , , �9  G� �9  H� ��  H� ��  G� �9  G�      C  , , �9  B� �9  C5 ��  C5 ��  B� �9  B�      C  , , �  G� �  H� �Y  H� �Y  G� �  G�      C  , , ��  G� ��  H� �m  H� �m  G� ��  G�      C  , , �  G� �  H� �Y  H� �Y  G� �  G�      C  , , �  B� �  C5 �Y  C5 �Y  B� �  B�      C  , , �  IW �  J �Y  J �Y  IW �  IW      C  , , �9  IW �9  J ��  J ��  IW �9  IW      C  , , �9  A# �9  A� ��  A� ��  A# �9  A#      C  , , ��  A# ��  A� �m  A� �m  A# ��  A#      C  , , �j  L �j  L� �  L� �  L �j  L      C  , , �  L �  L� �  L� �  L �  L      C  , , �%  B� �%  C5 ��  C5 ��  B� �%  B�      C  , , �%  A# �%  A� ��  A� ��  A# �%  A#      C  , , �~  L �~  L� �(  L� �(  L �~  L      C  , , �  IW �  J �Y  J �Y  IW �  IW      C  , , �  A# �  A� �Y  A� �Y  A# �  A#      C  , , ��  ;� ��  <- �~  <- �~  ;� ��  ;�      C  , , ��  IW ��  J �m  J �m  IW ��  IW      C  , , ��  L ��  L� �  L� �  L ��  L      C  , , �%  G� �%  H� ��  H� ��  G� �%  G�      C  , , ��  B� ��  C5 �m  C5 �m  B� ��  B�      C  , , ��  G� ��  H� �m  H� �m  G� ��  G�      C  , , �  A# �  A� �Y  A� �Y  A# �  A#      C  , , �%  IW �%  J ��  J ��  IW �%  IW      C  , , �9  G� �9  H� ��  H� ��  G� �9  G�      C  , , ��  IW ��  J �m  J �m  IW ��  IW      C  , , �9  %� �9  &a ��  &a ��  %� �9  %�      C  , , �  6 �  6� �Y  6� �Y  6 �  6      C  , , �  (� �  )1 �Y  )1 �Y  (� �  (�      C  , , �  +W �  , �Y  , �Y  +W �  +W      C  , , �9  (� �9  )1 ��  )1 ��  (� �9  (�      C  , , �  +W �  , �Y  , �Y  +W �  +W      C  , , �9  6 �9  6� ��  6� ��  6 �9  6      C  , , �9  )� �9  *� ��  *� ��  )� �9  )�      C  , , ��  ' ��  '� �m  '� �m  ' ��  '      C  , , �%  ' �%  '� ��  '� ��  ' �%  '      C  , , ��  ' ��  '� �m  '� �m  ' ��  '      C  , , �  4� �  5M �Y  5M �Y  4� �  4�      C  , , �   � �  !C �6  !C �6   � �   �      C  , , �9  +W �9  , ��  , ��  +W �9  +W      C  , , �%  )� �%  *� ��  *� ��  )� �%  )�      C  , , �9  4� �9  5M ��  5M ��  4� �9  4�      C  , , ��  )� ��  *� �m  *� �m  )� ��  )�      C  , , �$   � �$  !C ��  !C ��   � �$   �      C  , , ��   � ��  !C �l  !C �l   � ��   �      C  , , �  ' �  '� �Y  '� �Y  ' �  '      C  , , �  )� �  *� �Y  *� �Y  )� �  )�      C  , , �  3; �  3� �Y  3� �Y  3; �  3;      C  , , �9  %� �9  &a ��  &a ��  %� �9  %�      C  , , ��  (� ��  )1 �m  )1 �m  (� ��  (�      C  , , �  )� �  *� �Y  *� �Y  )� �  )�      C  , , �9  3; �9  3� ��  3� ��  3; �9  3;      C  , , �%  %� �%  &a ��  &a ��  %� �%  %�      C  , , ��  %� ��  &a �m  &a �m  %� ��  %�      C  , , �9  )� �9  *� ��  *� ��  )� �9  )�      C  , , �  1� �  2} �Y  2} �Y  1� �  1�      C  , , ��  )� ��  *� �m  *� �m  )� ��  )�      C  , , �%  +W �%  , ��  , ��  +W �%  +W      C  , , ��  +W ��  , �m  , �m  +W ��  +W      C  , , ��  %� ��  &a �m  &a �m  %� ��  %�      C  , , �  %� �  &a �Y  &a �Y  %� �  %�      C  , , �9  1� �9  2} ��  2} ��  1� �9  1�      C  , , �  (� �  )1 �Y  )1 �Y  (� �  (�      C  , , ��   � ��  !C �n  !C �n   � ��   �      C  , , �  0k �  1 �Y  1 �Y  0k �  0k      C  , , ��   � ��  !C �  !C �   � ��   �      C  , , �  %� �  &a �Y  &a �Y  %� �  %�      C  , , �9  (� �9  )1 ��  )1 ��  (� �9  (�      C  , , �9  0k �9  1 ��  1 ��  0k �9  0k      C  , , �%  (� �%  )1 ��  )1 ��  (� �%  (�      C  , , ��  (� ��  )1 �m  )1 �m  (� ��  (�      C  , , �9  ' �9  '� ��  '� ��  ' �9  '      C  , , �\   � �\  !C �  !C �   � �\   �      C  , , �  ' �  '� �Y  '� �Y  ' �  '      C  , , �9  +W �9  , ��  , ��  +W �9  +W      C  , , �j  #2 �j  #� �  #� �  #2 �j  #2      C  , , �9  ' �9  '� ��  '� ��  ' �9  '      C  , , �  #2 �  #� �  #� �  #2 �  #2      C  , , �~  #2 �~  #� �(  #� �(  #2 �~  #2      C  , , ��  #2 ��  #� �  #� �  #2 ��  #2      C  , , ��  +W ��  , �m  , �m  +W ��  +W      C  , , �   � �  !C �<  !C �<   � �   �      C  , , �M  )� �M  *� ��  *� ��  )� �M  )�      C  , , ��  )� ��  *� ��  *� ��  )� ��  )�      C  , , �M  ' �M  '� ��  '� ��  ' �M  '      C  , , �M  4� �M  5M ��  5M ��  4� �M  4�      C  , , ��  4� ��  5M ��  5M ��  4� ��  4�      C  , , ��  ' ��  '� ��  '� ��  ' ��  '      C  , , ��   � ��  !C �r  !C �r   � ��   �      C  , , ��  +W ��  , ��  , ��  +W ��  +W      C  , , �u  +W �u  , �  , �  +W �u  +W      C  , , ��  %� ��  &a ��  &a ��  %� ��  %�      C  , , �u  %� �u  &a �  &a �  %� �u  %�      C  , , ��  4� ��  5M ��  5M ��  4� ��  4�      C  , , �u  4� �u  5M �  5M �  4� �u  4�      C  , , �0   � �0  !C ��  !C ��   � �0   �      C  , , ��  %� ��  &a ��  &a ��  %� ��  %�      C  , , �  #2 �  #� �<  #� �<  #2 �  #2      C  , , �0  #2 �0  #� ��  #� ��  #2 �0  #2      C  , , �a  %� �a  &a �  &a �  %� �a  %�      C  , , �M  +W �M  , ��  , ��  +W �M  +W      C  , , �M  3; �M  3� ��  3� ��  3; �M  3;      C  , , ��  3; ��  3� ��  3� ��  3; ��  3;      C  , , �M  )� �M  *� ��  *� ��  )� �M  )�      C  , , ��  )� ��  *� ��  *� ��  )� ��  )�      C  , , ��  +W ��  , ��  , ��  +W ��  +W      C  , , �a  (� �a  )1 �  )1 �  (� �a  (�      C  , , �a  +W �a  , �  , �  +W �a  +W      C  , , �a  %� �a  &a �  &a �  %� �a  %�      C  , , ��  3; ��  3� ��  3� ��  3; ��  3;      C  , , �u  3; �u  3� �  3� �  3; �u  3;      C  , , ��  ' ��  '� ��  '� ��  ' ��  '      C  , , �M  %� �M  &a ��  &a ��  %� �M  %�      C  , , ��  %� ��  &a ��  &a ��  %� ��  %�      C  , , ��  )� ��  *� ��  *� ��  )� ��  )�      C  , , �u  )� �u  *� �  *� �  )� �u  )�      C  , , �u  ' �u  '� �  '� �  ' �u  '      C  , , �M  1� �M  2} ��  2} ��  1� �M  1�      C  , , ��  1� ��  2} ��  2} ��  1� ��  1�      C  , , ��  (� ��  )1 ��  )1 ��  (� ��  (�      C  , , �u  (� �u  )1 �  )1 �  (� �u  (�      C  , , ��  %� ��  &a ��  &a ��  %� ��  %�      C  , , �M  (� �M  )1 ��  )1 ��  (� �M  (�      C  , , ��  (� ��  )1 ��  )1 ��  (� ��  (�      C  , , �u  %� �u  &a �  &a �  %� �u  %�      C  , , ��  1� ��  2} ��  2} ��  1� ��  1�      C  , , �u  1� �u  2} �  2} �  1� �u  1�      C  , , �  #2 �  #� �P  #� �P  #2 �  #2      C  , , �M  (� �M  )1 ��  )1 ��  (� �M  (�      C  , , ��  (� ��  )1 ��  )1 ��  (� ��  (�      C  , , �M  %� �M  &a ��  &a ��  %� �M  %�      C  , , �b   � �b  !C �  !C �   � �b   �      C  , , �  #2 �  #� ��  #� ��  #2 �  #2      C  , , �M  0k �M  1 ��  1 ��  0k �M  0k      C  , , ��  0k ��  1 ��  1 ��  0k ��  0k      C  , , �    � �   !C ��  !C ��   � �    �      C  , , ��  #2 ��  #� �d  #� �d  #2 ��  #2      C  , , �a  )� �a  *� �  *� �  )� �a  )�      C  , , �a  )� �a  *� �  *� �  )� �a  )�      C  , , ��  (� ��  )1 ��  )1 ��  (� ��  (�      C  , , �a  ' �a  '� �  '� �  ' �a  '      C  , , ��  0k ��  1 ��  1 ��  0k ��  0k      C  , , �u  0k �u  1 �  1 �  0k �u  0k      C  , , �u  (� �u  )1 �  )1 �  (� �u  (�      C  , , �M  6 �M  6� ��  6� ��  6 �M  6      C  , , ��  6 ��  6� ��  6� ��  6 ��  6      C  , , ��  )� ��  *� ��  *� ��  )� ��  )�      C  , , �u  )� �u  *� �  *� �  )� �u  )�      C  , , ��   � ��  !C �  !C �   � ��   �      C  , , �a  ' �a  '� �  '� �  ' �a  '      C  , , �M  ' �M  '� ��  '� ��  ' �M  '      C  , , ��  ' ��  '� ��  '� ��  ' ��  '      C  , , �`   � �`  !C �
  !C �
   � �`   �      C  , , ��  +W ��  , ��  , ��  +W ��  +W      C  , , �u  +W �u  , �  , �  +W �u  +W      C  , , ��   � ��  !C �B  !C �B   � ��   �      C  , , �M  +W �M  , ��  , ��  +W �M  +W      C  , , �a  +W �a  , �  , �  +W �a  +W      C  , , ��  ' ��  '� ��  '� ��  ' ��  '      C  , , �u  ' �u  '� �  '� �  ' �u  '      C  , , ��  6 ��  6� ��  6� ��  6 ��  6      C  , , �u  6 �u  6� �  6� �  6 �u  6      C  , , ��  +W ��  , ��  , ��  +W ��  +W      C  , , �a  (� �a  )1 �  )1 �  (� �a  (�      C  , , 
�  >� 
�  ?> *  ?> *  >� 
�  >�      C  , , 	;  G� 	;  H� 	�  H� 	�  G� 	;  G�      C  , , �  G� �  H� �  H� �  G� �  G�      C  , , O  G� O  H� �  H� �  G� O  G�      C  , , �  IW �  J o  J o  IW �  IW      C  , , �  L �  L� �  L� �  L �  L      C  , , �  L �  L� >  L� >  L �  L      C  , , 
  L 
  L� �  L� �  L 
  L      C  , , �  A# �  A� o  A� o  A# �  A#      C  , , 	;  B� 	;  C5 	�  C5 	�  B� 	;  B�      C  , , 	;  IW 	;  J 	�  J 	�  IW 	;  IW      C  , , �  A# �  A� [  A� [  A# �  A#      C  , , O  A# O  A� �  A� �  A# O  A#      C  , , �  IW �  J [  J [  IW �  IW      C  , , �  IW �  J [  J [  IW �  IW      C  , , O  IW O  J �  J �  IW O  IW      C  , , O  IW O  J �  J �  IW O  IW      C  , , �  IW �  J o  J o  IW �  IW      C  , , �  B� �  C5 [  C5 [  B� �  B�      C  , , O  B� O  C5 �  C5 �  B� O  B�      C  , , �  B� �  C5 o  C5 o  B� �  B�      C  , , 	;  G� 	;  H� 	�  H� 	�  G� 	;  G�      C  , , 	;  IW 	;  J 	�  J 	�  IW 	;  IW      C  , , �  IW �  J �  J �  IW �  IW      C  , , �  G� �  H� o  H� o  G� �  G�      C  , , �  G� �  H� o  H� o  G� �  G�      C  , , L  ;� L  <- �  <- �  ;� L  ;�      C  , , �  ;� �  <- �  <- �  ;� �  ;�      C  , , �  G� �  H� [  H� [  G� �  G�      C  , , O  G� O  H� �  H� �  G� O  G�      C  , , �  B� �  C5 o  C5 o  B� �  B�      C  , , 	;  A# 	;  A� 	�  A� 	�  A# 	;  A#      C  , , 
�  L 
�  L� *  L� *  L 
�  L      C  , , �  A# �  A� o  A� o  A# �  A#      C  , , �  G� �  H� [  H� [  G� �  G�      C  , , �D  >� �D  ?> ��  ?> ��  >� �D  >�      C  , , ��  IW ��  J �3  J �3  IW ��  IW      C  , , '  IW '  J �  J �  IW '  IW      C  , , '  A# '  A� �  A� �  A# '  A#      C  , , �  B� �  C5 ��  C5 ��  B� �  B�      C  , , �  B� �  C5 G  C5 G  B� �  B�      C  , , ��  B� ��  C5 �3  C5 �3  B� ��  B�      C  , , ��  A# ��  A� ��  A� ��  A# ��  A#      C  , , ��  IW ��  J ��  J ��  IW ��  IW      C  , , �  IW �  J G  J G  IW �  IW      C  , , ��  G� ��  H� ��  H� ��  G� ��  G�      C  , , �  G� �  H� G  H� G  G� �  G�      C  , , �  A# �  A� ��  A� ��  A# �  A#      C  , , ��  IW ��  J ��  J ��  IW ��  IW      C  , , �  IW �  J G  J G  IW �  IW      C  , , ��  B� ��  C5 �3  C5 �3  B� ��  B�      C  , , '  B� '  C5 �  C5 �  B� '  B�      C  , , ��  G� ��  H� �3  H� �3  G� ��  G�      C  , , '  G� '  H� �  H� �  G� '  G�      C  , , '  B� '  C5 �  C5 �  B� '  B�      C  , , ��  ;� ��  <-  X  <-  X  ;� ��  ;�      C  , , ��  G� ��  H� �3  H� �3  G� ��  G�      C  , , '  G� '  H� �  H� �  G� '  G�      C  , ,  X  L  X  L�   L�   L  X  L      C  , , ��  B� ��  C5 ��  C5 ��  B� ��  B�      C  , , �  IW �  J ��  J ��  IW �  IW      C  , , �  G� �  H� ��  H� ��  G� �  G�      C  , , ��  A# ��  A� �3  A� �3  A# ��  A#      C  , , �  IW �  J ��  J ��  IW �  IW      C  , , �  A# �  A� G  A� G  A# �  A#      C  , , ��  L ��  L� �x  L� �x  L ��  L      C  , , ��  A# ��  A� �3  A� �3  A# ��  A#      C  , , �D  L �D  L� ��  L� ��  L �D  L      C  , , �  L �  L� �  L� �  L �  L      C  , , l  L l  L�   L�   L l  L      C  , , '  A# '  A� �  A� �  A# '  A#      C  , , ��  IW ��  J �3  J �3  IW ��  IW      C  , , �  G� �  H� ��  H� ��  G� �  G�      C  , , '  IW '  J �  J �  IW '  IW      C  , , ��  G� ��  H� ��  H� ��  G� ��  G�      C  , , �  G� �  H� G  H� G  G� �  G�      C  , , ��  )� ��  *� ��  *� ��  )� ��  )�      C  , , �  )� �  *� G  *� G  )� �  )�      C  , , �  (� �  )1 ��  )1 ��  (� �  (�      C  , , �  6 �  6� ��  6� ��  6 �  6      C  , , �  ' �  '� G  '� G  ' �  '      C  , , ��   � ��  !C ��  !C ��   � ��   �      C  , , �   � �  !C F  !C F   � �   �      C  , , �  +W �  , ��  , ��  +W �  +W      C  , , ��  4� ��  5M �3  5M �3  4� ��  4�      C  , , '  4� '  5M �  5M �  4� '  4�      C  , , �  +W �  , ��  , ��  +W �  +W      C  , , ��  ' ��  '� �3  '� �3  ' ��  '      C  , , '  ' '  '� �  '� �  ' '  '      C  , , ��  )� ��  *� �3  *� �3  )� ��  )�      C  , , ��   � ��  !C �x  !C �x   � ��   �      C  , , �  (� �  )1 ��  )1 ��  (� �  (�      C  , , �  4� �  5M ��  5M ��  4� �  4�      C  , , ��  ' ��  '� �3  '� �3  ' ��  '      C  , , '  ' '  '� �  '� �  ' '  '      C  , , l   � l  !C   !C    � l   �      C  , , �  ' �  '� ��  '� ��  ' �  '      C  , , '  )� '  *� �  *� �  )� '  )�      C  , , ��  3; ��  3� �3  3� �3  3; ��  3;      C  , , '  3; '  3� �  3� �  3; '  3;      C  , , �  )� �  *� G  *� G  )� �  )�      C  , , �6   � �6  !C ��  !C ��   � �6   �      C  , , ��  )� ��  *� �3  *� �3  )� ��  )�      C  , , ��  (� ��  )1 ��  )1 ��  (� ��  (�      C  , , �  (� �  )1 G  )1 G  (� �  (�      C  , , ��  %� ��  &a �3  &a �3  %� ��  %�      C  , , �  3; �  3� ��  3� ��  3; �  3;      C  , , '  %� '  &a �  &a �  %� '  %�      C  , , '  )� '  *� �  *� �  )� '  )�      C  , , ��  %� ��  &a ��  &a ��  %� ��  %�      C  , , �  %� �  &a G  &a G  %� �  %�      C  , , ��  +W ��  , ��  , ��  +W ��  +W      C  , , �  +W �  , G  , G  +W �  +W      C  , , ��  %� ��  &a ��  &a ��  %� ��  %�      C  , , ��  1� ��  2} �3  2} �3  1� ��  1�      C  , , '  1� '  2} �  2} �  1� '  1�      C  , , ��  +W ��  , �3  , �3  +W ��  +W      C  , , ��  (� ��  )1 �3  )1 �3  (� ��  (�      C  , , �  %� �  &a ��  &a ��  %� �  %�      C  , , �  ' �  '� ��  '� ��  ' �  '      C  , , �  1� �  2} ��  2} ��  1� �  1�      C  , , '  (� '  )1 �  )1 �  (� '  (�      C  , , ��  %� ��  &a �3  &a �3  %� ��  %�      C  , , '  %� '  &a �  &a �  %� '  %�      C  , , �  )� �  *� ��  *� ��  )� �  )�      C  , , '  +W '  , �  , �  +W '  +W      C  , , ��  #2 ��  #� �x  #� �x  #2 ��  #2      C  , , l  #2 l  #�   #�   #2 l  #2      C  , , ��  0k ��  1 �3  1 �3  0k ��  0k      C  , , '  0k '  1 �  1 �  0k '  0k      C  , , �f   � �f  !C �  !C �   � �f   �      C  , ,    �   !C �  !C �   �    �      C  , , ��  ' ��  '� ��  '� ��  ' ��  '      C  , , �  ' �  '� G  '� G  ' �  '      C  , , �  )� �  *� ��  *� ��  )� �  )�      C  , , �D  #2 �D  #� ��  #� ��  #2 �D  #2      C  , , �  0k �  1 ��  1 ��  0k �  0k      C  , , ��  +W ��  , ��  , ��  +W ��  +W      C  , , �  +W �  , G  , G  +W �  +W      C  , , �  #2 �  #� �  #� �  #2 �  #2      C  , , �  %� �  &a G  &a G  %� �  %�      C  , , ��  (� ��  )1 �3  )1 �3  (� ��  (�      C  , , '  (� '  )1 �  )1 �  (� '  (�      C  , , ��  )� ��  *� ��  *� ��  )� ��  )�      C  , ,  X  #2  X  #�   #�   #2  X  #2      C  , , �  %� �  &a ��  &a ��  %� �  %�      C  , , ��  +W ��  , �3  , �3  +W ��  +W      C  , , '  +W '  , �  , �  +W '  +W      C  , , ��  6 ��  6� �3  6� �3  6 ��  6      C  , , '  6 '  6� �  6� �  6 '  6      C  , ,  �   �  �  !C H  !C H   �  �   �      C  , , ��  (� ��  )1 ��  )1 ��  (� ��  (�      C  , , �  (� �  )1 G  )1 G  (� �  (�      C  , , ��  ' ��  '� ��  '� ��  ' ��  '      C  , , 	;  (� 	;  )1 	�  )1 	�  (� 	;  (�      C  , , �  (� �  )1 �  )1 �  (� �  (�      C  , , 	;  %� 	;  &a 	�  &a 	�  %� 	;  %�      C  , , �  +W �  , [  , [  +W �  +W      C  , , �  3; �  3� [  3� [  3; �  3;      C  , , O  3; O  3� �  3� �  3; O  3;      C  , , 	;  +W 	;  , 	�  , 	�  +W 	;  +W      C  , , �  %� �  &a o  &a o  %� �  %�      C  , , �  +W �  , �  , �  +W �  +W      C  , , <   � <  !C �  !C �   � <   �      C  , , �  +W �  , [  , [  +W �  +W      C  , , O  +W O  , �  , �  +W O  +W      C  , , �  (� �  )1 [  )1 [  (� �  (�      C  , , O  +W O  , �  , �  +W O  +W      C  , , �  6 �  6� [  6� [  6 �  6      C  , , O  6 O  6� �  6� �  6 O  6      C  , , �  1� �  2} o  2} o  1� �  1�      C  , , O  (� O  )1 �  )1 �  (� O  (�      C  , , 	;  )� 	;  *� 	�  *� 	�  )� 	;  )�      C  , , �  )� �  *� �  *� �  )� �  )�      C  , , �  %� �  &a [  &a [  %� �  %�      C  , , O  %� O  &a �  &a �  %� O  %�      C  , , �  (� �  )1 o  )1 o  (� �  (�      C  , , �  ' �  '� [  '� [  ' �  '      C  , , O  ' O  '� �  '� �  ' O  '      C  , , 	;  (� 	;  )1 	�  )1 	�  (� 	;  (�      C  , , �  1� �  2} [  2} [  1� �  1�      C  , , O  1� O  2} �  2} �  1� O  1�      C  , , �  %� �  &a o  &a o  %� �  %�      C  , , 
:   � 
:  !C 
�  !C 
�   � 
:   �      C  , , �  +W �  , o  , o  +W �  +W      C  , , �  )� �  *� [  *� [  )� �  )�      C  , , O  )� O  *� �  *� �  )� O  )�      C  , , �  4� �  5M o  5M o  4� �  4�      C  , , �   � �  !C �  !C �   � �   �      C  , , 
  #2 
  #� �  #� �  #2 
  #2      C  , , �  ' �  '� o  '� o  ' �  '      C  , , �  %� �  &a �  &a �  %� �  %�      C  , , �  0k �  1 o  1 o  0k �  0k      C  , , �  ' �  '� o  '� o  ' �  '      C  , , �   � �  !C L  !C L   � �   �      C  , , 
   � 
  !C �  !C �   � 
   �      C  , , 	;  )� 	;  *� 	�  *� 	�  )� 	;  )�      C  , , 	;  ' 	;  '� 	�  '� 	�  ' 	;  '      C  , , �  ' �  '� �  '� �  ' �  '      C  , , �  (� �  )1 [  )1 [  (� �  (�      C  , , �  #2 �  #� �  #� �  #2 �  #2      C  , , �  4� �  5M [  5M [  4� �  4�      C  , , �  0k �  1 [  1 [  0k �  0k      C  , , O  0k O  1 �  1 �  0k O  0k      C  , , O  4� O  5M �  5M �  4� O  4�      C  , , O  (� O  )1 �  )1 �  (� O  (�      C  , , 	;  +W 	;  , 	�  , 	�  +W 	;  +W      C  , , 
�  #2 
�  #� *  #� *  #2 
�  #2      C  , , �  )� �  *� [  *� [  )� �  )�      C  , , O  )� O  *� �  *� �  )� O  )�      C  , , �   � �  !C ~  !C ~   � �   �      C  , , �  ' �  '� [  '� [  ' �  '      C  , , O  ' O  '� �  '� �  ' O  '      C  , , r   � r  !C   !C    � r   �      C  , , �  %� �  &a [  &a [  %� �  %�      C  , , �  #2 �  #� >  #� >  #2 �  #2      C  , , �  (� �  )1 o  )1 o  (� �  (�      C  , , �  +W �  , o  , o  +W �  +W      C  , , O  %� O  &a �  &a �  %� O  %�      C  , , �  3; �  3� o  3� o  3; �  3;      C  , , �  )� �  *� o  *� o  )� �  )�      C  , , �  )� �  *� o  *� o  )� �  )�      C  , , 	;  ' 	;  '� 	�  '� 	�  ' 	;  '      C  , , 	;  %� 	;  &a 	�  &a 	�  %� 	;  %�      C  , , �  6 �  6� o  6� o  6 �  6      ^   , �c  M� �c  P7 ��  P7 ��  M� �c  M�      ^   , ��  M� ��  P7 �]  P7 �]  M� ��  M�      ^   , ~  V� ~  X� (  X� (  V� ~  V�      ^   , y  e� y  n� a  n� a  e� y  e�      ^   , �  e� �  n� �  n� �  e� �  e�      ^   , ;  e� ;  n� #  n� #  e� ;  e�      ^   , 
�  e� 
�  n� �  n� �  e� 
�  e�      ^   , �  M� �  P7 �3  P7 �3  M� �  M�      ^   , �9  M� �9  P7 ��  P7 ��  M� �9  M�      ^   , ��  M� ��  P7 o  P7 o  M� ��  M�      ^   , ��  M� ��  P7 �  P7 �  M� ��  M�      ^   , �  M� �  P7 �3  P7 �3  M� �  M�      ^   , �9  M� �9  P7 ��  P7 ��  M� �9  M�      ^   , ��  M� ��  P7 o  P7 o  M� ��  M�      ^   , u  M� u  P7 
  P7 
  M� u  M�      ^   , 	  M� 	  P7 �  P7 �  M� 	  M�      ^   , u  M� u  P7 
  P7 
  M� u  M�      ^   , ��  M� ��  P7 �  P7 �  M� ��  M�      ^   , �  p� �  ym �  ym �  p� �  p�      ^   , �  p� �  ym �S  ym �S  p� �  p�      ^   , �A  p� �A  ym ��  ym ��  p� �A  p�      ^   , �{  $w �{  -A �+  -A �+  $w �{  $w      ^   , �  $w �  -A ��  -A ��  $w �  $w      ^   , ��  $w ��  -A �g  -A �g  $w ��  $w      ^   , �U  $w �U  -A   -A   $w �U  $w      ^   , �  $w �  -A 
�  -A 
�  $w �  $w      ^   , �  $w �  -A A  -A A  $w �  $w      ^   ,  �  p�  �  ym �  ym �  p�  �  p�      ^   , �g  p� �g  ym �  ym �  p� �g  p�      ^   , �  p� �  ym �?  ym �?  p� �  p�      ^   , �-  p� �-  ym ��  ym ��  p� �-  p�      ^   , ��  p� ��  ym  {  ym  {  p� ��  p�      ^   , ��  $w ��  -A �  -A �  $w ��  $w      ^   , �  $w �  -A �?  -A �?  $w �  $w      ^   , �-  $w �-  -A ��  -A ��  $w �-  $w      ^   , ��  $w ��  -A  {  -A  {  $w ��  $w      ^   , i  $w i  -A   -A   $w i  $w      ^   ,   $w   -A �  -A �  $w   $w      ^   , i  p� i  ym   ym   p� i  p�      ^   , ��  p� ��  ym �  ym �  p� ��  p�      ^   , �  p� �  ym ��  ym ��  p� �  p�      ^   , ��  p� ��  ym �g  ym �g  p� ��  p�      ^   , �U  p� �U  ym   ym   p� �U  p�      ^   , �g  $w �g  -A �  -A �  $w �g  $w      ^   , �  $w �  -A �  -A �  $w �  $w      ^   , �  $w �  -A �S  -A �S  $w �  $w      ^   , �A  $w �A  -A ��  -A ��  $w �A  $w      ^   ,  �  $w  �  -A �  -A �  $w  �  $w      ^   , }  $w }  -A -  -A -  $w }  $w      ^   , �  p� �  ym 
�  ym 
�  p� �  p�      ^   , �{  p� �{  ym �+  ym �+  p� �{  p�      ^   , �  e� �  n� �?  n� �?  e� �  e�      ^   , �-  e� �-  n� ��  n� ��  e� �-  e�      ^   , ��  e� ��  n�  {  n�  {  e� ��  e�      ^   , ��  /+ ��  7� �  7� �  /+ ��  /+      ^   , �  /+ �  7� �?  7� �?  /+ �  /+      ^   , �-  /+ �-  7� ��  7� ��  /+ �-  /+      ^   , ��  /+ ��  7�  {  7�  {  /+ ��  /+      ^   , i  /+ i  7�   7�   /+ i  /+      ^   ,   /+   7� �  7� �  /+   /+      ^   , i  e� i  n�   n�   e� i  e�      ^   , ��  e� ��  n� �  n� �  e� ��  e�      ^   , ��  p� ��  ym �  ym �  p� ��  p�   	   B   !     ^  ��  e� ��  ^t   	   B   !     ^  ��  e� ��  ^t   	   B   !     ^  �#  e� �#  ^t   	   B   !     ^  �I  8@ �I  ?p   	   B   !     ^  ��  8@ ��  ?p   	   B   !     ^  ��  8@ ��  ?p   	   B   !     ^  �#  8@ �#  ?p   	   B   !     ^  �  8@ �  ?p   	   B   !     ^  _  8@ _  ?p   	   B   !     ^  �  e� �  ^t   	   B   !     ^  �I  e� �I  ^t   	   B   !     @  �  b �  b   	   B   !     @  �J  b �4  b   	   B   !     @  ��  b ��  b   	   B   !     @  �  ;� �  ;�   	   B   !     @  �"  ;� �8  ;�   	   B   !     @  ��  ;� ��  ;�   	   B   !     @  �^  ;� �t  ;�   	   B   !     @  �  ;�   ;�   	   B   !     @  �  ;� �  ;�   	   B   !     @  �  b p  b   	   B   !     @  �  b ��  b   	   B   !     ^  ��  C� ��  HS   	   B   !     ^  7  C� 7  HS   	   B   !     ^  �5  S\ �5  P�   	   B   !     ^  ��  ZU ��  U�   	   B   !     ^  �  ZU �  U�   	   B   !     ^  K  ZU K  U�   	   B   !      �  �  ]� �  e�   	   B   !      �  �  ]� �  fq   	   B   !      �  /  ^ /  f   	   B   !      �  m  ]� m  f!   	   B   !      �  �  l� �  o�   	   B   !      �  m  l� m  o�   	   B   !      �  �  l� �  o�      B   , �`  P� �`  R0 ��  R0 ��  P� �`  P�      B   , �`  R0 �`  W� ��  W� ��  R0 �`  R0      B   , �`  y� �`  { ��  { ��  y� �`  y�      B   , �`  pX �`  y� ��  y� ��  pX �`  pX      B   , �`  X� �`  ^t ��  ^t ��  X� �`  X�      B   , �`  $, �`  -� ��  -� ��  $, �`  $,      B   , �`  K� �`  L� ��  L� ��  K� �`  K�      B   , �`  "� �`  $, ��  $, ��  "� �`  "�      B   , �`  F< �`  K� ��  K� ��  F< �`  F<      B   , �  X� �  ^t <  ^t <  X� �  X�      B   , "  X� "  ^t �  ^t �  X� "  X�      B   , �  X� �  ^t z  ^t z  X� �  X�      B   , �t  X� �t  ^t ��  ^t ��  X� �t  X�      B   ,   X�   ^t p  ^t p  X�   X�      B   , ��  al ��  b� ��  b� ��  al ��  al      B   , <  al <  b� �  b� �  al <  al      B   , �t  P� �t  R0 ��  R0 ��  P� �t  P�      B   ,   P�   R0 p  R0 p  P�   P�      B   , �t  R0 �t  W� ��  W� ��  R0 �t  R0      B   ,   R0   W� p  W� p  R0   R0      B   , ��  P� ��  R0 �H  R0 �H  P� ��  P�      B   , �  P� �  R0 �  R0 �  P� �  P�      B   , ��  R0 ��  W� �H  W� �H  R0 ��  R0      B   , �  R0 �  W� �  W� �  R0 �  R0      B   , ��  P� ��  R0 \  R0 \  P� ��  P�      B   , �  P� �  R0 �  R0 �  P� �  P�      B   , ��  R0 ��  W� \  W� \  R0 ��  R0      B   , �  R0 �  W� �  W� �  R0 �  R0      B   , ��  y� ��  { �H  { �H  y� ��  y�      B   , �  y� �  { �  { �  y� �  y�      B   , ��  pX ��  y� �H  y� �H  pX ��  pX      B   , �  pX �  y� �  y� �  pX �  pX      B   , �t  y� �t  { ��  { ��  y� �t  y�      B   ,   y�   { p  { p  y�   y�      B   , �t  pX �t  y� ��  y� ��  pX �t  pX      B   ,   pX   y� p  y� p  pX   pX      B   , ��  y� ��  { \  { \  y� ��  y�      B   , �  y� �  { �  { �  y� �  y�      B   , ��  pX ��  y� \  y� \  pX ��  pX      B   , �  pX �  y� �  y� �  pX �  pX      B   , �t  e� �t  o ��  o ��  e� �t  e�      B   ,   e�   o p  o p  e�   e�      B   , �  X� �  ^t �  ^t �  X� �  X�      B   , ��  ^t ��  _� \  _� \  ^t ��  ^t      B   , "  e� "  o �  o �  e� "  e�      B   , �  e� �  o <  o <  e� �  e�      B   , �  e� �  o z  o z  e� �  e�      B   , `  e� `  o �  o �  e� `  e�      B   , ��  X� ��  ^t \  ^t \  X� ��  X�      B   , �  a� �  b� 7  b� 7  a� �  a�      B   , �  n} �  o� �  o� �  n} �  n}      B   , `  X� `  ^t �  ^t �  X� `  X�      B   , ��  R0 ��  W� �   W� �   R0 ��  R0      B   , �<  P� �<  R0 �  R0 �  P� �<  P�      B   , ��  P� ��  R0 �4  R0 �4  P� ��  P�      B   , ��  X� ��  ^t �4  ^t �4  X� ��  X�      B   , �$  R0 �$  W� �  W� �  R0 �$  R0      B   , �  y� �  { �  { �  y� �  y�      B   , �L  y� �L  { ��  { ��  y� �L  y�      B   , �  pX �  y� ��  y� ��  pX �  pX      B   , �  P� �  R0 ��  R0 ��  P� �  P�      B   , �  y� �  { �n  { �n  y� �  y�      B   , �  pX �  y� �  y� �  pX �  pX      B   , �L  pX �L  y� ��  y� ��  pX �L  pX      B   , �8  R0 �8  W� �  W� �  R0 �8  R0      B   , ��  R0 ��  W� �4  W� �4  R0 ��  R0      B   , �  pX �  y� �n  y� �n  pX �  pX      B   , �8  y� �8  { �  { �  y� �8  y�      B   , ��  y� ��  { �4  { �4  y� ��  y�      B   , ��  X� ��  ^t �   ^t �   X� ��  X�      B   , �  X� �  ^t ��  ^t ��  X� �  X�      B   , �  y� �  { ��  { ��  y� �  y�      B   , �8  pX �8  y� �  y� �  pX �8  pX      B   , ��  pX ��  y� �4  y� �4  pX ��  pX      B   , �  R0 �  W� ��  W� ��  R0 �  R0      B   , �  P� �  R0 �  R0 �  P� �  P�      B   , �  pX �  y� ��  y� ��  pX �  pX      B   , ��  y� ��  { �   { �   y� ��  y�      B   , �8  X� �8  ^t �  ^t �  X� �8  X�      B   , �L  P� �L  R0 ��  R0 ��  P� �L  P�      B   , �b  al �b  b� �  b� �  al �b  al      B   , �$  y� �$  { �  { �  y� �$  y�      B   , ��  pX ��  y� �   y� �   pX ��  pX      B   , �  R0 �  W� �n  W� �n  R0 �  R0      B   , �   al �   b� �J  b� �J  al �   al      B   , �  P� �  R0 �n  R0 �n  P� �  P�      B   , �$  pX �$  y� �  y� �  pX �$  pX      B   , �8  e� �8  o �  o �  e� �8  e�      B   , ��  e� ��  o �4  o �4  e� ��  e�      B   , �  R0 �  W� �  W� �  R0 �  R0      B   , �L  R0 �L  W� ��  W� ��  R0 �L  R0      B   , �  e� �  o ��  o ��  e� �  e�      B   , �  y� �  { ��  { ��  y� �  y�      B   , ��  P� ��  R0 �   R0 �   P� ��  P�      B   , �  R0 �  W� ��  W� ��  R0 �  R0      B   , �$  X� �$  ^t �  ^t �  X� �$  X�      B   , ��  ^t ��  _� �   _� �   ^t ��  ^t      B   , ��  al ��  b� �  b� �  al ��  al      B   , �8  P� �8  R0 �  R0 �  P� �8  P�      B   , �$  P� �$  R0 �  R0 �  P� �$  P�      B   , �  F< �  K� ��  K� ��  F< �  F<      B   , �8  F< �8  K� �  K� �  F< �8  F<      B   , ��  F< ��  K� �4  K� �4  F< ��  F<      B   , �  ?p �  D� ��  D� ��  ?p �  ?p      B   , �  "� �  $, ��  $, ��  "� �  "�      B   , �8  "� �8  $, �  $, �  "� �8  "�      B   , ��  "� ��  $, �4  $, �4  "� ��  "�      B   , �  K� �  L� �n  L� �n  K� �  K�      B   , �  K� �  L� �  L� �  K� �  K�      B   , �L  K� �L  L� ��  L� ��  K� �L  K�      B   , �8  ?p �8  D� �  D� �  ?p �8  ?p      B   , ��  ?p ��  D� �4  D� �4  ?p ��  ?p      B   , �  $, �  -� ��  -� ��  $, �  $,      B   , �8  $, �8  -� �  -� �  $, �8  $,      B   , ��  $, ��  -� �4  -� �4  $, ��  $,      B   , �  K� �  L� ��  L� ��  K� �  K�      B   , �8  K� �8  L� �  L� �  K� �8  K�      B   , �$  K� �$  L� �  L� �  K� �$  K�      B   , �  F< �  K� �n  K� �n  F< �  F<      B   , �  F< �  K� �  K� �  F< �  F<      B   , �  "� �  $, �n  $, �n  "� �  "�      B   , �  "� �  $, �  $, �  "� �  "�      B   , �L  "� �L  $, ��  $, ��  "� �L  "�      B   , �L  F< �L  K� ��  K� ��  F< �L  F<      B   , ��  K� ��  L� �   L� �   K� ��  K�      B   , �  >b �  ?p �  ?p �  >b �  >b      B   , ��  K� ��  L� �4  L� �4  K� ��  K�      B   , �  ;8 �  <x ��  <x ��  ;8 �  ;8      B   , �  $, �  -� �n  -� �n  $, �  $,      B   , �  $, �  -� �  -� �  $, �  $,      B   , �L  $, �L  -� ��  -� ��  $, �L  $,      B   , �"  ;8 �"  <x �l  <x �l  ;8 �"  ;8      B   , �$  "� �$  $, �  $, �  "� �$  "�      B   , ��  "� ��  $, �   $, �   "� ��  "�      B   , �  >b �  ?p �n  ?p �n  >b �  >b      B   , ��  ;8 ��  <x �
  <x �
  ;8 ��  ;8      B   , �  .� �  8@ ��  8@ ��  .� �  .�      B   , �8  .� �8  8@ �  8@ �  .� �8  .�      B   , ��  .� ��  8@ �4  8@ �4  .� ��  .�      B   , �  ?p �  D� �  D� �  ?p �  ?p      B   , �$  F< �$  K� �  K� �  F< �$  F<      B   , �L  ?p �L  D� ��  D� ��  ?p �L  ?p      B   , ��  F< ��  K� �   K� �   F< ��  F<      B   , �  ?p �  D� �n  D� �n  ?p �  ?p      B   , �$  $, �$  -� �  -� �  $, �$  $,      B   , ��  $, ��  -� �   -� �   $, ��  $,      B   , ��  >b ��  ?p �H  ?p �H  >b ��  >b      B   , 
&  >b 
&  ?p �  ?p �  >b 
&  >b      B   , �  F< �  K� �  K� �  F< �  F<      B   , :  F< :  K� �  K� �  F< :  F<      B   , �  K� �  L�   L�   K� �  K�      B   ,   ?p   D� p  D� p  ?p   ?p      B   , �t  $, �t  -� ��  -� ��  $, �t  $,      B   ,   $,   -� p  -� p  $,   $,      B   , �  $, �  -�   -�   $, �  $,      B   , �  ?p �  D�   D�   ?p �  ?p      B   , 
&  ?p 
&  D� �  D� �  ?p 
&  ?p      B   , ��  "� ��  $, \  $, \  "� ��  "�      B   , �  "� �  $, �  $, �  "� �  "�      B   , :  "� :  $, �  $, �  "� :  "�      B   , ��  ?p ��  D� �H  D� �H  ?p ��  ?p      B   , �t  ?p �t  D� ��  D� ��  ?p �t  ?p      B   , ��  K� ��  L� \  L� \  K� ��  K�      B   , ��  "� ��  $, �H  $, �H  "� ��  "�      B   , �  "� �  $, �  $, �  "� �  "�      B   , 
&  "� 
&  $, �  $, �  "� 
&  "�      B   , �  K� �  L� �  L� �  K� �  K�      B   , ��  K� ��  L� �H  L� �H  K� ��  K�      B   , �  K� �  L� �  L� �  K� �  K�      B   , 
&  K� 
&  L� �  L� �  K� 
&  K�      B   , :  K� :  L� �  L� �  K� :  K�      B   , ��  $, ��  -� \  -� \  $, ��  $,      B   , �  $, �  -� �  -� �  $, �  $,      B   , :  $, :  -� �  -� �  $, :  $,      B   , ��  $, ��  -� �H  -� �H  $, ��  $,      B   , �  $, �  -� �  -� �  $, �  $,      B   , 
&  $, 
&  -� �  -� �  $, 
&  $,      B   , �^  ;8 �^  <x  �  <x  �  ;8 �^  ;8      B   , �  ;8 �  <x F  <x F  ;8 �  ;8      B   , �  ;8 �  <x �  <x �  ;8 �  ;8      B   , �t  F< �t  K� ��  K� ��  F< �t  F<      B   ,   F<   K� p  K� p  F<   F<      B   , �  F< �  K�   K�   F< �  F<      B   , �t  K� �t  L� ��  L� ��  K� �t  K�      B   , ��  F< ��  K� �H  K� �H  F< ��  F<      B   , �t  .� �t  8@ ��  8@ ��  .� �t  .�      B   ,   .�   8@ p  8@ p  .�   .�      B   , �  .� �  8@   8@   .� �  .�      B   , �t  "� �t  $, ��  $, ��  "� �t  "�      B   ,   "�   $, p  $, p  "�   "�      B   , �  "� �  $,   $,   "� �  "�      B   , �  F< �  K� �  K� �  F< �  F<      B   , 
&  F< 
&  K� �  K� �  F< 
&  F<      B   , �  ?p �  D� �  D� �  ?p �  ?p      B   ,   K�   L� p  L� p  K�   K�      B   , ��  F< ��  K� \  K� \  F< ��  F<      A   , �4  Y� �4  ]� ��  ]� ��  Y� �4  Y�      A   , ��  @8 ��  D  �t  D  �t  @8 ��  @8      A   , ��  R� ��  V� �t  V� �t  R� ��  R�      A   , �4  G �4  J� ��  J� ��  G �4  G      A   , �4  R� �4  V� ��  V� ��  R� �4  R�      A   , ��  G ��  J� �t  J� �t  G ��  G      A   , ��  q  ��  x� �t  x� �t  q  ��  q       A   , �4  $� �4  ,� ��  ,� ��  $� �4  $�      A   , �4  q  �4  x� ��  x� ��  q  �4  q       A   , ��  $� ��  ,� �t  ,� �t  $� ��  $�      A   , �H  R� �H  V� ��  V� ��  R� �H  R�      A   , �  R� �  V� �  V� �  R� �  R�      A   , �  fl �  n< �  n< �  fl �  fl      A   , z  fl z  n< h  n< h  fl z  fl      A   , \  R� \  V�   V�   R� \  R�      A   , �  fl �  n< �  n< �  fl �  fl      A   , ��  R� ��  V� �  V� �  R� ��  R�      A   , 4  fl 4  n< "  n< "  fl 4  fl      A   , p  R� p  V� 
&  V� 
&  R� p  R�      A   , ��  Y� ��  ]� �  ]� �  Y� ��  Y�      A   , p  Y� p  ]� 
&  ]� 
&  Y� p  Y�      A   , \  q  \  x�   x�   q  \  q       A   , �H  q  �H  x� ��  x� ��  q  �H  q       A   , �  q  �  x� �  x� �  q  �  q       A   , �H  Y� �H  ]� ��  ]� ��  Y� �H  Y�      A   , ��  q  ��  x� �  x� �  q  ��  q       A   , �  Y� �  ]� �  ]� �  Y� �  Y�      A   , p  q  p  x� 
&  x� 
&  q  p  q       A   , �H  fl �H  n< ��  n< ��  fl �H  fl      A   , �  fl �  n< �  n< �  fl �  fl      A   , 4  Y� 4  ]� "  ]� "  Y� 4  Y�      A   , z  Y� z  ]� h  ]� h  Y� z  Y�      A   , �  Y� �  ]� �  ]� �  Y� �  Y�      A   , �  Y� �  ]� �  ]� �  Y� �  Y�      A   , �  q  �  x� �8  x� �8  q  �  q       A   , �   q  �   x� ��  x� ��  q  �   q       A   , ��  Y� ��  ]� �  ]� �  Y� ��  Y�      A   , �Z  q  �Z  x� �  x� �  q  �Z  q       A   , �n  R� �n  V� �$  V� �$  R� �n  R�      A   , ��  q  ��  x� �  x� �  q  ��  q       A   , �  q  �  x� ��  x� ��  q  �  q       A   , ��  q  ��  x� �`  x� �`  q  ��  q       A   , �  R� �  V� �8  V� �8  R� �  R�      A   , �   R� �   V� ��  V� ��  R� �   R�      A   , �n  q  �n  x� �$  x� �$  q  �n  q       A   , �  q  �  x� �L  x� �L  q  �  q       A   , �  Y� �  ]� ��  ]� ��  Y� �  Y�      A   , ��  Y� ��  ]� �`  ]� �`  Y� ��  Y�      A   , �Z  R� �Z  V� �  V� �  R� �Z  R�      A   , ��  R� ��  V� �  V� �  R� ��  R�      A   , ��  q  ��  x� �  x� �  q  ��  q       A   , �  fl �  n< ��  n< ��  fl �  fl      A   , ��  fl ��  n< �`  n< �`  fl ��  fl      A   , �  R� �  V� �L  V� �L  R� �  R�      A   , �  Y� �  ]� �L  ]� �L  Y� �  Y�      A   , �n  fl �n  n< �$  n< �$  fl �n  fl      A   , �n  Y� �n  ]� �$  ]� �$  Y� �n  Y�      A   , �  R� �  V� ��  V� ��  R� �  R�      A   , ��  R� ��  V� �`  V� �`  R� ��  R�      A   , ��  R� ��  V� �  V� �  R� ��  R�      A   , ��  $� ��  ,� �`  ,� �`  $� ��  $�      A   , �   G �   J� ��  J� ��  G �   G      A   , �  @8 �  D  ��  D  ��  @8 �  @8      A   , ��  @8 ��  D  �`  D  �`  @8 ��  @8      A   , ��  G ��  J� �  J� �  G ��  G      A   , �  G �  J� �L  J� �L  G �  G      A   , ��  $� ��  ,� �  ,� �  $� ��  $�      A   , �  $� �  ,� �8  ,� �8  $� �  $�      A   , �   $� �   ,� ��  ,� ��  $� �   $�      A   , �n  G �n  J� �$  J� �$  G �n  G      A   , �  G �  J� ��  J� ��  G �  G      A   , ��  $� ��  ,� �  ,� �  $� ��  $�      A   , �  $� �  ,� �L  ,� �L  $� �  $�      A   , ��  G ��  J� �`  J� �`  G ��  G      A   , �  @8 �  D  �8  D  �8  @8 �  @8      A   , �n  /� �n  7x �$  7x �$  /� �n  /�      A   , �  /� �  7x ��  7x ��  /� �  /�      A   , ��  /� ��  7x �`  7x �`  /� ��  /�      A   , �   @8 �   D  ��  D  ��  @8 �   @8      A   , �n  @8 �n  D  �$  D  �$  @8 �n  @8      A   , ��  @8 ��  D  �  D  �  @8 ��  @8      A   , ��  G ��  J� �  J� �  G ��  G      A   , �  G �  J� �8  J� �8  G �  G      A   , �n  $� �n  ,� �$  ,� �$  $� �n  $�      A   , �  $� �  ,� ��  ,� ��  $� �  $�      A   , ��  $� ��  ,� �  ,� �  $� ��  $�      A   , p  $� p  ,� 
&  ,� 
&  $� p  $�      A   ,   $�   ,� �  ,� �  $�   $�      A   , �  G �  J� �  J� �  G �  G      A   , \  $� \  ,�   ,�   $� \  $�      A   , �  $� �  ,� �  ,� �  $� �  $�      A   , �  G �  J� :  J� :  G �  G      A   , ��  G ��  J� �  J� �  G ��  G      A   , \  G \  J�   J�   G \  G      A   , �  G �  J� �  J� �  G �  G      A   , p  G p  J� 
&  J� 
&  G p  G      A   ,   G   J� �  J� �  G   G      A   , �  @8 �  D  �  D  �  @8 �  @8      A   , �H  $� �H  ,� ��  ,� ��  $� �H  $�      A   , �H  /� �H  7x ��  7x ��  /� �H  /�      A   , �  /� �  7x �  7x �  /� �  /�      A   , �  /� �  7x :  7x :  /� �  /�      A   , �  $� �  ,� �  ,� �  $� �  $�      A   , �  $� �  ,� :  ,� :  $� �  $�      A   , �  @8 �  D  :  D  :  @8 �  @8      A   , �  @8 �  D  �  D  �  @8 �  @8      A   , \  @8 \  D    D    @8 \  @8      A   , �H  @8 �H  D  ��  D  ��  @8 �H  @8      A   , �H  G �H  J� ��  J� ��  G �H  G      _   , ��  ^B ��  _� �  _� �  ^B ��  ^B      _   , �  ^B �  _� �R  _� �R  ^B �  ^B      _   , ��  >0 ��  ?� �  ?� �  >0 ��  >0      _   , �|  >0 �|  ?� �>  ?� �>  >0 �|  >0      _   , ��  >0 ��  ?� �z  ?� �z  >0 ��  >0      _   , 	�  >0 	�  ?� �  ?� �  >0 	�  >0      _   , �
  P� �
  Rb �  Rb �  P� �
  P�      _   , �|  y� �|  { ��  { ��  y� �|  y�      _   , �  aS �  b� i  b� i  aS �  aS      _   , h  nK h  o� �  o� �  nK h  nK      _   , �0  a: �0  b� ��  b� ��  a: �0  a:      _   , ��  a: ��  b� �|  b� �|  a: ��  a:      _   , �l  a: �l  b� �  b� �  a: �l  a:      _   , �R  ; �R  <� �   <� �   ; �R  ;      _   , ��  ; ��  <� �  <� �  ; ��  ;      _   , ��  ; ��  <� �<  <� �<  ; ��  ;      _   , �,  ; �,  <�  �  <�  �  ; �,  ;      _   , �  ; �  <� x  <� x  ; �  ;      _   , h  ; h  <�   <�   ; h  ;      _   , 
  a: 
  b� �  b� �  a: 
  a:      _   , �  a: �  b� �@  b� �@  a: �  a:      _   , �.  P� �.  R: �  R: �  P� �.  P�      _   , ��  P� ��  R: �>  R: �>  P� ��  P�      _   , �j  P� �j  R: ��  R: ��  P� �j  P�      _   , �  K� �  M �  M �  K� �  K�      _   , �.  K� �.  M �  M �  K� �.  K�      _   , ��  K� ��  M �>  M �>  K� ��  K�      _   , �j  K� �j  M ��  M ��  K� �j  K�      _   ,   K�   M z  M z  K�   K�      _   , �  K� �  M   M   K� �  K�      _   ,   P�   R: z  R: z  P�   P�      _   , �  P� �  R: �  R: �  P� �  P�      _   , �  P� �  R: �  R: �  P� �  P�      _   , �B  P� �B  R: ��  R: ��  P� �B  P�      _   , ��  P� ��  R: �R  R: �R  P� ��  P�      _   , �  K� �  M �  M �  K� �  K�      _   , �  K� �  M �*  M �*  K� �  K�      _   , �V  K� �V  M ��  M ��  K� �V  K�      _   , ��  K� ��  M f  M f  K� ��  K�      _   , �  K� �  M 	  M 	  K� �  K�      _   , 0  K� 0  M �  M �  K� 0  K�      _   , ~  P� ~  R: �  R: �  P� ~  P�      _   , �  P� �  R: �x  R: �x  P� �  P�      _   , �  P� �  R: �*  R: �*  P� �  P�      _   , �V  P� �V  R: ��  R: ��  P� �V  P�      _   , ��  P� ��  R: f  R: f  P� ��  P�      _   , �  K� �  M �x  M �x  K� �  K�      _   , �  K� �  M �  M �  K� �  K�      _   , �B  K� �B  M ��  M ��  K� �B  K�      _   , ��  K� ��  M �R  M �R  K� ��  K�      _   , ~  K� ~  M �  M �  K� ~  K�      _   , 
  K� 
  M �  M �  K� 
  K�      _   , �  P� �  R: 	  R: 	  P� �  P�      _   , �  P� �  R: �  R: �  P� �  P�      _   , �  y� �  { �  { �  y� �  y�      _   , �B  y� �B  { ��  { ��  y� �B  y�      _   , ��  y� ��  { �R  { �R  y� ��  y�      _   , �  "� �  $6 �  $6 �  "� �  "�      _   , �  "� �  $6 �*  $6 �*  "� �  "�      _   , �V  "� �V  $6 ��  $6 ��  "� �V  "�      _   , ��  "� ��  $6 f  $6 f  "� ��  "�      _   , �  "� �  $6 	  $6 	  "� �  "�      _   , 0  "� 0  $6 �  $6 �  "� 0  "�      _   , ~  y� ~  { �  { �  y� ~  y�      _   , �  y� �  { �x  { �x  y� �  y�      _   , �.  y� �.  { �  { �  y� �.  y�      _   , ��  y� ��  { �>  { �>  y� ��  y�      _   , �j  y� �j  { ��  { ��  y� �j  y�      _   , �  "� �  $6 �  $6 �  "� �  "�      _   , �.  "� �.  $6 �  $6 �  "� �.  "�      _   , ��  "� ��  $6 �>  $6 �>  "� ��  "�      _   , �j  "� �j  $6 ��  $6 ��  "� �j  "�      _   ,   "�   $6 z  $6 z  "�   "�      _   , �  "� �  $6   $6   "� �  "�      _   ,   y�   { z  { z  y�   y�      _   , �  y� �  { �  { �  y� �  y�      _   , �  y� �  { �*  { �*  y� �  y�      _   , �V  y� �V  { ��  { ��  y� �V  y�      _   , ��  y� ��  { f  { f  y� ��  y�      _   , �  "� �  $6 �x  $6 �x  "� �  "�      _   , �  "� �  $6 �  $6 �  "� �  "�      _   , �B  "� �B  $6 ��  $6 ��  "� �B  "�      _   , ��  "� ��  $6 �R  $6 �R  "� ��  "�      _   , ~  "� ~  $6 �  $6 �  "� ~  "�      _   , 
  "� 
  $6 �  $6 �  "� 
  "�      _   , �  y� �  { 	  { 	  y� �  y�      _   , �  y� �  { �  { �  y� �  y�      }  , , ��  Y ��  ^` �r  ^` �r  Y ��  Y      }  , , ��  FP ��  K� �r  K� �r  FP ��  FP      }  , , ��  RD ��  W� �r  W� �r  RD ��  RD      }  , , ��  $@ ��  -x �r  -x �r  $@ ��  $@      }  , , ��  pl ��  y� �r  y� �r  pl ��  pl      }  , , ��  RD ��  W� ��  W� ��  RD ��  RD      }  , , ^  RD ^  W� $  W� $  RD ^  RD      }  , , �6  RD �6  W� ��  W� ��  RD �6  RD      }  , , �  Y �  ^` 	�  ^` 	�  Y �  Y      }  , , �  RD �  W� �  W� �  RD �  RD      }  , , �J  Y �J  ^`   ^`   Y �J  Y      }  , , �J  RD �J  W�   W�   RD �J  RD      }  , , �  RD �  W� 	�  W� 	�  RD �  RD      }  , , �6  pl �6  y� ��  y� ��  pl �6  pl      }  , , ��  Y ��  ^` ��  ^` ��  Y ��  Y      }  , , �  pl �  y� �  y� �  pl �  pl      }  , , ��  pl ��  y� ��  y� ��  pl ��  pl      }  , , ^  pl ^  y� $  y� $  pl ^  pl      }  , , ^  Y ^  ^` $  ^` $  Y ^  Y      }  , , �J  pl �J  y�   y�   pl �J  pl      }  , , �  pl �  y� 	�  y� 	�  pl �  pl      }  , , ��  e� ��  n� ��  n� ��  e� ��  e�      }  , , ^  e� ^  n� $  n� $  e� ^  e�      }  , , �  RD �  W� ��  W� ��  RD �  RD      }  , , �  Y �  ^` ��  ^` ��  Y �  Y      }  , , ��  Y ��  ^` �  ^` �  Y ��  Y      }  , , �  RD �  W� �J  W� �J  RD �  RD      }  , , �p  RD �p  W� �6  W� �6  RD �p  RD      }  , , ��  pl ��  y� ��  y� ��  pl ��  pl      }  , , �  pl �  y� �^  y� �^  pl �  pl      }  , , �"  RD �"  W� ��  W� ��  RD �"  RD      }  , , �p  Y �p  ^` �6  ^` �6  Y �p  Y      }  , , ��  pl ��  y� �  y� �  pl ��  pl      }  , , �\  pl �\  y� �"  y� �"  pl �\  pl      }  , , �  pl �  y� �J  y� �J  pl �  pl      }  , , �"  pl �"  y� ��  y� ��  pl �"  pl      }  , , ��  RD ��  W� �  W� �  RD ��  RD      }  , , ��  RD ��  W� ��  W� ��  RD ��  RD      }  , , ��  pl ��  y� �  y� �  pl ��  pl      }  , , �  pl �  y� ��  y� ��  pl �  pl      }  , , �  RD �  W� �^  W� �^  RD �  RD      }  , , �  Y �  ^` �J  ^` �J  Y �  Y      }  , , �"  Y �"  ^` ��  ^` ��  Y �"  Y      }  , , �p  pl �p  y� �6  y� �6  pl �p  pl      }  , , �  e� �  n� �J  n� �J  e� �  e�      }  , , �"  e� �"  n� ��  n� ��  e� �"  e�      }  , , ��  RD ��  W� �  W� �  RD ��  RD      }  , , �\  RD �\  W� �"  W� �"  RD �\  RD      }  , , ��  e� ��  n� �  n� �  e� ��  e�      }  , , �  FP �  K� �J  K� �J  FP �  FP      }  , , �"  FP �"  K� ��  K� ��  FP �"  FP      }  , , �"  ?� �"  D� ��  D� ��  ?� �"  ?�      }  , , �  ?� �  D� �^  D� �^  ?� �  ?�      }  , , ��  $@ ��  -x �  -x �  $@ ��  $@      }  , , �  $@ �  -x �J  -x �J  $@ �  $@      }  , , �"  $@ �"  -x ��  -x ��  $@ �"  $@      }  , , �\  FP �\  K� �"  K� �"  FP �\  FP      }  , , ��  FP ��  K� ��  K� ��  FP ��  FP      }  , , �  FP �  K� �^  K� �^  FP �  FP      }  , , ��  ?� ��  D� ��  D� ��  ?� ��  ?�      }  , , �\  ?� �\  D� �"  D� �"  ?� �\  ?�      }  , , �\  $@ �\  -x �"  -x �"  $@ �\  $@      }  , , ��  $@ ��  -x ��  -x ��  $@ ��  $@      }  , , �  $@ �  -x �^  -x �^  $@ �  $@      }  , , ��  ?� ��  D� �  D� �  ?� ��  ?�      }  , , �p  FP �p  K� �6  K� �6  FP �p  FP      }  , , �  FP �  K� ��  K� ��  FP �  FP      }  , , �p  $@ �p  -x �6  -x �6  $@ �p  $@      }  , , �  $@ �  -x ��  -x ��  $@ �  $@      }  , , ��  .� ��  8, �  8, �  .� ��  .�      }  , , �  .� �  8, �J  8, �J  .� �  .�      }  , , �"  .� �"  8, ��  8, ��  .� �"  .�      }  , , �  ?� �  D� �J  D� �J  ?� �  ?�      }  , , ��  FP ��  K� �  K� �  FP ��  FP      }  , , ��  $@ ��  -x ��  -x ��  $@ ��  $@      }  , , ^  $@ ^  -x $  -x $  $@ ^  $@      }  , , �  $@ �  -x �  -x �  $@ �  $@      }  , , �J  FP �J  K�   K�   FP �J  FP      }  , , �  FP �  K� 	�  K� 	�  FP �  FP      }  , , �  FP �  K� L  K� L  FP �  FP      }  , , �  FP �  K� �  K� �  FP �  FP      }  , , �  ?� �  D� �  D� �  ?� �  ?�      }  , , ��  ?� ��  D� ��  D� ��  ?� ��  ?�      }  , , ^  ?� ^  D� $  D� $  ?� ^  ?�      }  , , �J  $@ �J  -x   -x   $@ �J  $@      }  , , �6  $@ �6  -x ��  -x ��  $@ �6  $@      }  , , �  $@ �  -x �  -x �  $@ �  $@      }  , , 	r  $@ 	r  -x 8  -x 8  $@ 	r  $@      }  , , �  $@ �  -x 	�  -x 	�  $@ �  $@      }  , , �  $@ �  -x L  -x L  $@ �  $@      }  , , �  ?� �  D� �  D� �  ?� �  ?�      }  , , �6  ?� �6  D� ��  D� ��  ?� �6  ?�      }  , , 	r  ?� 	r  D� 8  D� 8  ?� 	r  ?�      }  , , ��  FP ��  K� ��  K� ��  FP ��  FP      }  , , �6  FP �6  K� ��  K� ��  FP �6  FP      }  , , �  FP �  K� �  K� �  FP �  FP      }  , , ��  .� ��  8, ��  8, ��  .� ��  .�      }  , , ^  .� ^  8, $  8, $  .� ^  .�      }  , , �  .� �  8, �  8, �  .� �  .�      }  , , 	r  FP 	r  K� 8  K� 8  FP 	r  FP      }  , , ^  FP ^  K� $  K� $  FP ^  FP      D      �  eO out       D      �M  ^� vrst      D      �  |� vdd       D      ��  N� vss       D      �  N� vss       D      ��  |� vdd       D      �  b out       D      ��  b out       D      W  b out       D        B�        �  ;� out       D        B�        �  ;� out       D        B�        �Q  ;� out       D        B�        ��  ;� out       D        B�        �  ;� out       D        B�        
+  ;� out       D      �  b out       D      �}  b out       D      �  |� vdd       D      �"  |� vdd       D      �  |� vdd       D        B�        �   � vdd       D        B�        �J   � vdd       D        B�        ��   � vdd       D        B�        ��   � vdd       D        B�        $   � vdd       D        B�        	�   � vdd       D      	^  |� vdd       D      ��  |� vdd       D      �\  N� vss       D      ��  N� vss       D      �  N� vss       D        B�        ��  N� vss       D        B�        �r  N� vss       D        B�        �  N� vss       D        B�        ��  N� vss       D        B�        L  N� vss       D        B�        	�  N� vss       D      	6  N� vss       D      �  N� vss       D      �J  b in      D      ��  b in      D      ��  b in      D        B�        ��  ;� in      D        B�        �  ;� in      D        B�        �"  ;� in      D        B�        �  ;� in      D        B�        	^  ;� in      D        B�        �  ;� in      D      $  b in      D      �  b in      F      ��  n� 
vctrp       F      ��  LY 
vctrn       F      ��  T� vss       F      ��  Q� 
vctrn       F      ��  u vdd       F      �S  u vdd       F      ��  u vdd       F      ��  u vdd       F        B�        ��  (� vdd       F        B�        �{  (� vdd       F        B�        �  (� vdd       F        B�         �  (� vdd       F        B�        U  (� vdd       F        B�        �  (� vdd       F      -  u vdd       F      �  u vdd       F      �  z] 
vctrp       F      �O  z] 
vctrp       F      ��  z] 
vctrp       F        B�        �  #� 
vctrp       F        B�        �  #� 
vctrp       F        B�        ��  #� 
vctrp       F        B�        �Y  #� 
vctrp       F        B�        �  #� 
vctrp       F        B�        �  #� 
vctrp       F      �  z] 
vctrp       F      �  z] 
vctrp       F      ��  T� vss       F      �s  T� vss       F      �  T� vss       F        B�        �[  H� vss       F        B�        ��  H� vss       F        B�        ��  H� vss       F        B�         5  H� vss       F        B�        �  H� vss       F        B�        q  H� vss       F      �  T� vss       F      �7  T� vss       F      �  Q� 
vctrn       F      �@  Q� 
vctrn       F      ��  Q� 
vctrn       F        B�        �  LY 
vctrn       F        B�        �,  LY 
vctrn       F        B�        ��  LY 
vctrn       F        B�        �h  LY 
vctrn       F        B�          LY 
vctrn       F        B�        �  LY 
vctrn       F      |  Q� 
vctrn       F      �  Q� 
vctrn       D      �  e� out       D      �  ^� vrst      D      �E  |� vdd       D      �i  N� vss       D      �J  a� in      D      ��  a� in      D      ��  a� in      D        B�        ��  ;� in      D        B�        �  ;� in      D        B�        �"  ;� in      D        B�        �  ;� in      D        B�        	^  ;� in      D        B�        �  ;� in      D      $  a� in      D      �  a� in      D      �  a� out       D      ��  a� out       D      W  a� out       D        B�        �  ;� out       D        B�        �  ;� out       D        B�        �Q  ;� out       D        B�        ��  ;� out       D        B�        �  ;� out       D        B�        
+  ;� out       D      �  a� out       D      �}  a� out       D      �.  |� vdd       D      ��  |� vdd       D      �j  |� vdd       D        B�        �   � vdd       D        B�        �   � vdd       D        B�        �>   � vdd       D        B�        ��   � vdd       D        B�        z   � vdd       D        B�           � vdd       D        |� vdd       D      �  |� vdd       D      �  N� vss       D      �0  N� vss       D      ��  N� vss       D        B�        �  N� vss       D        B�        �<  N� vss       D        B�        ��  N� vss       D        B�        �x  N� vss       D        B�          N� vss       D        B�        �  N� vss       D      l  N� vss       D      ��  N� vss       F   , ֛  P� ֛  R0 �"  R0 �"  P� ֛  P�      F   , �a  S\ �a  T� �u  T� �u  S\ �a  S\      F      �>  LY 
vctrn       F      ��  T� vss       F      �>  Q� 
vctrn       F      �  u vdd       F      ��  Q� 
vctrn       F      �  T� vss       F      �f  z� 
vctrp       F      �  z� 
vctrp       F      �  z� 
vctrp       F        B�        ��  #Z 
vctrp       F        B�        �h  #Z 
vctrp       F        B�        �  #Z 
vctrp       F        B�        ��  #Z 
vctrp       F        B�        B  #Z 
vctrp       F        B�        	�  #Z 
vctrp       F      	@  z� 
vctrp       F      ��  z� 
vctrp       F      �k  Q� 
vctrn       F      �	  Q� 
vctrn       F      �  Q� 
vctrn       F        B�        ��  LY 
vctrn       F        B�        �c  LY 
vctrn       F        B�        �  LY 
vctrn       F        B�        ��  LY 
vctrn       F        B�        =  LY 
vctrn       F        B�        	�  LY 
vctrn       F      	E  Q� 
vctrn       F      ��  Q� 
vctrn       F      �>  T� vss       F      ��  T� vss       F      z  T� vss       F        B�        ��  H� vss       F        B�        �  H� vss       F        B�        �.  H� vss       F        B�        ��  H� vss       F        B�        j  H� vss       F        B�        
  H� vss       F      	  T� vss       F      �  T� vss       