VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_Onchip_RCO
  CLASS BLOCK ;
  FOREIGN tt_um_Onchip_RCO ;
  ORIGIN 203.340 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT -59.510 224.760 -59.210 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT -56.750 224.760 -56.450 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT -62.270 224.760 -61.970 225.760 ;
    END
  END rst_n
  PIN ua[0]
    PORT
      LAYER met4 ;
        RECT -51.530 0.000 -50.630 1.000 ;
    END
  END ua[0]
  PIN ua[2]
    PORT
      LAYER met4 ;
        RECT -90.170 0.000 -89.270 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    PORT
      LAYER met4 ;
        RECT -109.490 0.000 -108.590 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    PORT
      LAYER met4 ;
        RECT -128.810 0.000 -127.910 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT -148.130 0.000 -147.230 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT -167.450 0.000 -166.550 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT -186.770 0.000 -185.870 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 2.100000 ;
    PORT
      LAYER met4 ;
        RECT -65.030 224.760 -64.730 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT -67.790 224.760 -67.490 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    PORT
      LAYER met4 ;
        RECT -70.550 224.760 -70.250 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    PORT
      LAYER met4 ;
        RECT -73.310 224.760 -73.010 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    PORT
      LAYER met4 ;
        RECT -76.070 224.760 -75.770 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    PORT
      LAYER met4 ;
        RECT -78.830 224.760 -78.530 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    PORT
      LAYER met4 ;
        RECT -81.590 224.760 -81.290 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    PORT
      LAYER met4 ;
        RECT -84.350 224.760 -84.050 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    PORT
      LAYER met4 ;
        RECT -87.110 224.760 -86.810 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    PORT
      LAYER met4 ;
        RECT -89.870 224.760 -89.570 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    PORT
      LAYER met4 ;
        RECT -92.630 224.760 -92.330 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    PORT
      LAYER met4 ;
        RECT -95.390 224.760 -95.090 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    PORT
      LAYER met4 ;
        RECT -98.150 224.760 -97.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    PORT
      LAYER met4 ;
        RECT -100.910 224.760 -100.610 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    PORT
      LAYER met4 ;
        RECT -103.670 224.760 -103.370 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    PORT
      LAYER met4 ;
        RECT -106.430 224.760 -106.130 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -153.350 224.760 -153.050 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -156.110 224.760 -155.810 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -158.870 224.760 -158.570 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -161.630 224.760 -161.330 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -164.390 224.760 -164.090 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -167.150 224.760 -166.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -169.910 224.760 -169.610 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -172.670 224.760 -172.370 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -131.270 224.760 -130.970 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -134.030 224.760 -133.730 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -136.790 224.760 -136.490 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -139.550 224.760 -139.250 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -142.310 224.760 -142.010 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -145.070 224.760 -144.770 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -147.830 224.760 -147.530 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -150.590 224.760 -150.290 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -109.190 224.760 -108.890 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -111.950 224.760 -111.650 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -114.710 224.760 -114.410 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -117.470 224.760 -117.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -120.230 224.760 -119.930 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -122.990 224.760 -122.690 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -125.750 224.760 -125.450 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNAGATEAREA 9.450000 ;
    ANTENNADIFFAREA 16.455999 ;
    PORT
      LAYER met4 ;
        RECT -128.510 224.760 -128.210 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNAGATEAREA 15.400000 ;
    ANTENNADIFFAREA 24.855999 ;
    PORT
      LAYER met4 ;
        RECT -202.340 5.000 -200.340 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -199.340 5.000 -197.340 220.760 ;
    END
  END VGND
  PIN ua[1]
    ANTENNADIFFAREA 1.800000 ;
    PORT
      LAYER met4 ;
        RECT -70.850 0.000 -69.950 1.000 ;
    END
  END ua[1]
  OBS
      LAYER nwell ;
        RECT -180.910 8.050 -66.995 189.485 ;
      LAYER li1 ;
        RECT -180.600 8.230 -67.365 189.175 ;
      LAYER met1 ;
        RECT -187.450 8.230 -64.580 194.195 ;
      LAYER met2 ;
        RECT -187.450 8.230 -64.580 194.195 ;
      LAYER met3 ;
        RECT -202.340 8.230 -62.195 194.195 ;
      LAYER met4 ;
        RECT -197.340 224.360 -173.070 224.760 ;
        RECT -171.970 224.360 -170.310 224.760 ;
        RECT -169.210 224.360 -167.550 224.760 ;
        RECT -166.450 224.360 -164.790 224.760 ;
        RECT -163.690 224.360 -162.030 224.760 ;
        RECT -160.930 224.360 -159.270 224.760 ;
        RECT -158.170 224.360 -156.510 224.760 ;
        RECT -155.410 224.360 -153.750 224.760 ;
        RECT -152.650 224.360 -150.990 224.760 ;
        RECT -149.890 224.360 -148.230 224.760 ;
        RECT -147.130 224.360 -145.470 224.760 ;
        RECT -144.370 224.360 -142.710 224.760 ;
        RECT -141.610 224.360 -139.950 224.760 ;
        RECT -138.850 224.360 -137.190 224.760 ;
        RECT -136.090 224.360 -134.430 224.760 ;
        RECT -133.330 224.360 -131.670 224.760 ;
        RECT -130.570 224.360 -128.910 224.760 ;
        RECT -127.810 224.360 -126.150 224.760 ;
        RECT -125.050 224.360 -123.390 224.760 ;
        RECT -122.290 224.360 -120.630 224.760 ;
        RECT -119.530 224.360 -117.870 224.760 ;
        RECT -116.770 224.360 -115.110 224.760 ;
        RECT -114.010 224.360 -112.350 224.760 ;
        RECT -111.250 224.360 -109.590 224.760 ;
        RECT -108.490 224.360 -106.830 224.760 ;
        RECT -105.730 224.360 -104.070 224.760 ;
        RECT -102.970 224.360 -101.310 224.760 ;
        RECT -100.210 224.360 -98.550 224.760 ;
        RECT -97.450 224.360 -95.790 224.760 ;
        RECT -94.690 224.360 -93.030 224.760 ;
        RECT -91.930 224.360 -90.270 224.760 ;
        RECT -89.170 224.360 -87.510 224.760 ;
        RECT -86.410 224.360 -84.750 224.760 ;
        RECT -83.650 224.360 -81.990 224.760 ;
        RECT -80.890 224.360 -79.230 224.760 ;
        RECT -78.130 224.360 -76.470 224.760 ;
        RECT -75.370 224.360 -73.710 224.760 ;
        RECT -72.610 224.360 -70.950 224.760 ;
        RECT -69.850 224.360 -68.190 224.760 ;
        RECT -67.090 224.360 -65.430 224.760 ;
        RECT -64.330 224.360 -62.670 224.760 ;
        RECT -61.570 224.360 -59.910 224.760 ;
        RECT -58.810 224.360 -57.150 224.760 ;
        RECT -56.050 224.360 -50.625 224.760 ;
        RECT -197.340 221.160 -50.625 224.360 ;
        RECT -196.940 4.600 -50.625 221.160 ;
        RECT -197.340 1.400 -50.625 4.600 ;
        RECT -197.340 0.000 -187.170 1.400 ;
        RECT -185.470 0.000 -167.850 1.400 ;
        RECT -166.150 0.000 -148.530 1.400 ;
        RECT -146.830 0.000 -129.210 1.400 ;
        RECT -127.510 0.000 -109.890 1.400 ;
        RECT -108.190 0.000 -90.570 1.400 ;
        RECT -88.870 0.000 -71.250 1.400 ;
        RECT -69.550 0.000 -51.930 1.400 ;
  END
END tt_um_Onchip_RCO
END LIBRARY

