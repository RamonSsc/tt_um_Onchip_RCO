magic
tech sky130a
timestamp 1762644065
<< checkpaint >>
<< end >>
