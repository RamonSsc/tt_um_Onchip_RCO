magic
tech sky130a
timestamp 1762644065
<< checkpaint >>
rect 0 0 1 2
<< l70d20 >>
rect 0 0 1 2
<< l71d20 >>
rect 0 0 1 2
<< end >>
